// Copyright (C) 2017  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 17.1.1 Internal Build 593 12/11/2017 SJ Lite Edition"

// DATE "03/06/2018 12:30:33"

// 
// Device: Altera 5CSEMA4U23C6 Package UFBGA672
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module spw_babasu (
	autostart_external_connection_export,
	clk_clk,
	currentstate_external_connection_export,
	data_i_external_connection_export,
	data_o_external_connection_export,
	flags_external_connection_export,
	link_disable_external_connection_export,
	link_start_external_connection_export,
	pll_0_locked_export,
	pll_0_outclk0_clk,
	rd_data_external_connection_export,
	reset_reset_n,
	rx_empty_external_connection_export,
	spill_enable_external_connection_export,
	tick_in_external_connection_export,
	tick_out_external_connection_export,
	time_in_external_connection_export,
	time_out_external_connection_export,
	tx_clk_div_external_connection_export,
	tx_full_external_connection_export,
	wr_data_external_connection_export)/* synthesis synthesis_greybox=0 */;
output 	autostart_external_connection_export;
input 	clk_clk;
input 	[2:0] currentstate_external_connection_export;
output 	[8:0] data_i_external_connection_export;
input 	[8:0] data_o_external_connection_export;
input 	[10:0] flags_external_connection_export;
output 	link_disable_external_connection_export;
output 	link_start_external_connection_export;
output 	pll_0_locked_export;
output 	pll_0_outclk0_clk;
output 	rd_data_external_connection_export;
input 	reset_reset_n;
input 	rx_empty_external_connection_export;
output 	spill_enable_external_connection_export;
output 	tick_in_external_connection_export;
input 	tick_out_external_connection_export;
output 	[7:0] time_in_external_connection_export;
input 	[7:0] time_out_external_connection_export;
output 	[6:0] tx_clk_div_external_connection_export;
input 	tx_full_external_connection_export;
output 	wr_data_external_connection_export;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \hps_0|fpga_interfaces|h2f_rst_n[0] ;
wire \hps_0|fpga_interfaces|h2f_ARVALID[0] ;
wire \hps_0|fpga_interfaces|h2f_AWVALID[0] ;
wire \hps_0|fpga_interfaces|h2f_BREADY[0] ;
wire \hps_0|fpga_interfaces|h2f_RREADY[0] ;
wire \hps_0|fpga_interfaces|h2f_WLAST[0] ;
wire \hps_0|fpga_interfaces|h2f_WVALID[0] ;
wire \hps_0|fpga_interfaces|h2f_ARADDR[0] ;
wire \hps_0|fpga_interfaces|h2f_ARADDR[1] ;
wire \hps_0|fpga_interfaces|h2f_ARADDR[2] ;
wire \hps_0|fpga_interfaces|h2f_ARADDR[3] ;
wire \hps_0|fpga_interfaces|h2f_ARADDR[4] ;
wire \hps_0|fpga_interfaces|h2f_ARADDR[5] ;
wire \hps_0|fpga_interfaces|h2f_ARADDR[6] ;
wire \hps_0|fpga_interfaces|h2f_ARADDR[7] ;
wire \hps_0|fpga_interfaces|h2f_ARADDR[8] ;
wire \hps_0|fpga_interfaces|h2f_ARBURST[0] ;
wire \hps_0|fpga_interfaces|h2f_ARBURST[1] ;
wire \hps_0|fpga_interfaces|h2f_ARID[0] ;
wire \hps_0|fpga_interfaces|h2f_ARID[1] ;
wire \hps_0|fpga_interfaces|h2f_ARID[2] ;
wire \hps_0|fpga_interfaces|h2f_ARID[3] ;
wire \hps_0|fpga_interfaces|h2f_ARID[4] ;
wire \hps_0|fpga_interfaces|h2f_ARID[5] ;
wire \hps_0|fpga_interfaces|h2f_ARID[6] ;
wire \hps_0|fpga_interfaces|h2f_ARID[7] ;
wire \hps_0|fpga_interfaces|h2f_ARID[8] ;
wire \hps_0|fpga_interfaces|h2f_ARID[9] ;
wire \hps_0|fpga_interfaces|h2f_ARID[10] ;
wire \hps_0|fpga_interfaces|h2f_ARID[11] ;
wire \hps_0|fpga_interfaces|h2f_ARLEN[0] ;
wire \hps_0|fpga_interfaces|h2f_ARLEN[1] ;
wire \hps_0|fpga_interfaces|h2f_ARLEN[2] ;
wire \hps_0|fpga_interfaces|h2f_ARLEN[3] ;
wire \hps_0|fpga_interfaces|h2f_ARSIZE[0] ;
wire \hps_0|fpga_interfaces|h2f_ARSIZE[1] ;
wire \hps_0|fpga_interfaces|h2f_ARSIZE[2] ;
wire \hps_0|fpga_interfaces|h2f_AWADDR[0] ;
wire \hps_0|fpga_interfaces|h2f_AWADDR[1] ;
wire \hps_0|fpga_interfaces|h2f_AWADDR[2] ;
wire \hps_0|fpga_interfaces|h2f_AWADDR[3] ;
wire \hps_0|fpga_interfaces|h2f_AWADDR[4] ;
wire \hps_0|fpga_interfaces|h2f_AWADDR[5] ;
wire \hps_0|fpga_interfaces|h2f_AWADDR[6] ;
wire \hps_0|fpga_interfaces|h2f_AWADDR[7] ;
wire \hps_0|fpga_interfaces|h2f_AWADDR[8] ;
wire \hps_0|fpga_interfaces|h2f_AWBURST[0] ;
wire \hps_0|fpga_interfaces|h2f_AWBURST[1] ;
wire \hps_0|fpga_interfaces|h2f_AWID[0] ;
wire \hps_0|fpga_interfaces|h2f_AWID[1] ;
wire \hps_0|fpga_interfaces|h2f_AWID[2] ;
wire \hps_0|fpga_interfaces|h2f_AWID[3] ;
wire \hps_0|fpga_interfaces|h2f_AWID[4] ;
wire \hps_0|fpga_interfaces|h2f_AWID[5] ;
wire \hps_0|fpga_interfaces|h2f_AWID[6] ;
wire \hps_0|fpga_interfaces|h2f_AWID[7] ;
wire \hps_0|fpga_interfaces|h2f_AWID[8] ;
wire \hps_0|fpga_interfaces|h2f_AWID[9] ;
wire \hps_0|fpga_interfaces|h2f_AWID[10] ;
wire \hps_0|fpga_interfaces|h2f_AWID[11] ;
wire \hps_0|fpga_interfaces|h2f_AWLEN[0] ;
wire \hps_0|fpga_interfaces|h2f_AWLEN[1] ;
wire \hps_0|fpga_interfaces|h2f_AWLEN[2] ;
wire \hps_0|fpga_interfaces|h2f_AWLEN[3] ;
wire \hps_0|fpga_interfaces|h2f_AWSIZE[0] ;
wire \hps_0|fpga_interfaces|h2f_AWSIZE[1] ;
wire \hps_0|fpga_interfaces|h2f_AWSIZE[2] ;
wire \hps_0|fpga_interfaces|h2f_WDATA[0] ;
wire \hps_0|fpga_interfaces|h2f_WDATA[1] ;
wire \hps_0|fpga_interfaces|h2f_WDATA[2] ;
wire \hps_0|fpga_interfaces|h2f_WDATA[3] ;
wire \hps_0|fpga_interfaces|h2f_WDATA[4] ;
wire \hps_0|fpga_interfaces|h2f_WDATA[5] ;
wire \hps_0|fpga_interfaces|h2f_WDATA[6] ;
wire \hps_0|fpga_interfaces|h2f_WDATA[7] ;
wire \hps_0|fpga_interfaces|h2f_WDATA[8] ;
wire \hps_0|fpga_interfaces|h2f_WSTRB[0] ;
wire \hps_0|fpga_interfaces|h2f_WSTRB[1] ;
wire \hps_0|fpga_interfaces|h2f_WSTRB[2] ;
wire \hps_0|fpga_interfaces|h2f_WSTRB[3] ;
wire \pll_0|altera_pll_i|outclk_wire[0] ;
wire \pll_0|altera_pll_i|locked_wire[0] ;
wire \autostart|data_out~q ;
wire \data_i|data_out[0]~q ;
wire \data_i|data_out[1]~q ;
wire \data_i|data_out[2]~q ;
wire \data_i|data_out[3]~q ;
wire \data_i|data_out[4]~q ;
wire \data_i|data_out[5]~q ;
wire \data_i|data_out[6]~q ;
wire \data_i|data_out[7]~q ;
wire \data_i|data_out[8]~q ;
wire \link_disable|data_out~q ;
wire \link_start|data_out~q ;
wire \rd_data|data_out~q ;
wire \spill_enable|data_out~q ;
wire \tick_in|data_out~q ;
wire \time_in|data_out[0]~q ;
wire \time_in|data_out[1]~q ;
wire \time_in|data_out[2]~q ;
wire \time_in|data_out[3]~q ;
wire \time_in|data_out[4]~q ;
wire \time_in|data_out[5]~q ;
wire \time_in|data_out[6]~q ;
wire \time_in|data_out[7]~q ;
wire \tx_clk_div|data_out[0]~q ;
wire \tx_clk_div|data_out[1]~q ;
wire \tx_clk_div|data_out[2]~q ;
wire \tx_clk_div|data_out[3]~q ;
wire \tx_clk_div|data_out[4]~q ;
wire \tx_clk_div|data_out[5]~q ;
wire \tx_clk_div|data_out[6]~q ;
wire \wr_data|data_out~q ;
wire \mm_interconnect_0|link_disable_s1_translator|wait_latency_counter[1]~q ;
wire \mm_interconnect_0|link_disable_s1_translator|wait_latency_counter[0]~q ;
wire \mm_interconnect_0|tx_clk_div_s1_translator|wait_latency_counter[1]~q ;
wire \mm_interconnect_0|tx_clk_div_s1_translator|wait_latency_counter[0]~q ;
wire \mm_interconnect_0|spill_enable_s1_translator|wait_latency_counter[1]~q ;
wire \mm_interconnect_0|spill_enable_s1_translator|wait_latency_counter[0]~q ;
wire \mm_interconnect_0|tick_in_s1_translator|wait_latency_counter[1]~q ;
wire \mm_interconnect_0|tick_in_s1_translator|wait_latency_counter[0]~q ;
wire \mm_interconnect_0|time_in_s1_translator|wait_latency_counter[1]~q ;
wire \mm_interconnect_0|time_in_s1_translator|wait_latency_counter[0]~q ;
wire \mm_interconnect_0|data_i_s1_translator|wait_latency_counter[1]~q ;
wire \mm_interconnect_0|data_i_s1_translator|wait_latency_counter[0]~q ;
wire \mm_interconnect_0|rd_data_s1_translator|wait_latency_counter[1]~q ;
wire \mm_interconnect_0|rd_data_s1_translator|wait_latency_counter[0]~q ;
wire \mm_interconnect_0|link_start_s1_translator|wait_latency_counter[1]~q ;
wire \mm_interconnect_0|link_start_s1_translator|wait_latency_counter[0]~q ;
wire \mm_interconnect_0|autostart_s1_translator|wait_latency_counter[1]~q ;
wire \mm_interconnect_0|autostart_s1_translator|wait_latency_counter[0]~q ;
wire \mm_interconnect_0|wr_data_s1_translator|wait_latency_counter[1]~q ;
wire \mm_interconnect_0|wr_data_s1_translator|wait_latency_counter[0]~q ;
wire \mm_interconnect_0|hps_0_h2f_axi_master_rd_limiter|cmd_sink_ready~0_combout ;
wire \mm_interconnect_0|hps_0_h2f_axi_master_wr_limiter|nonposted_cmd_accepted~0_combout ;
wire \mm_interconnect_0|rsp_mux|WideOr1~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload[0]~combout ;
wire \mm_interconnect_0|rsp_mux_001|WideOr1~combout ;
wire \mm_interconnect_0|hps_0_h2f_axi_master_wr_limiter|nonposted_cmd_accepted~1_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[105]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[106]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[107]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[108]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[109]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[110]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[111]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[112]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[113]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[114]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[115]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[116]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[0]~20_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~30_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~38_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~45_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~52_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~59_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~66_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~72_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~75_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~76_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~77_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[105]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[106]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[107]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[108]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[109]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[110]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[111]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[112]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[113]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[114]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[115]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[116]~combout ;
wire \mm_interconnect_0|autostart_s1_agent|m0_write~combout ;
wire \mm_interconnect_0|autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ;
wire \mm_interconnect_0|autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ;
wire \mm_interconnect_0|autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ;
wire \rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \mm_interconnect_0|data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ;
wire \mm_interconnect_0|data_i_s1_agent|m0_write~combout ;
wire \mm_interconnect_0|data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ;
wire \mm_interconnect_0|data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ;
wire \mm_interconnect_0|data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[1]~q ;
wire \mm_interconnect_0|data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[2]~q ;
wire \mm_interconnect_0|data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[3]~q ;
wire \mm_interconnect_0|data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[4]~q ;
wire \mm_interconnect_0|data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[5]~q ;
wire \mm_interconnect_0|data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[6]~q ;
wire \mm_interconnect_0|data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[7]~q ;
wire \mm_interconnect_0|data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[8]~q ;
wire \mm_interconnect_0|link_disable_s1_agent|m0_write~combout ;
wire \mm_interconnect_0|link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ;
wire \mm_interconnect_0|link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ;
wire \mm_interconnect_0|link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ;
wire \mm_interconnect_0|link_start_s1_agent|m0_write~combout ;
wire \mm_interconnect_0|link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ;
wire \mm_interconnect_0|link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ;
wire \mm_interconnect_0|link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ;
wire \mm_interconnect_0|rd_data_s1_agent|m0_write~combout ;
wire \mm_interconnect_0|rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ;
wire \mm_interconnect_0|rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ;
wire \mm_interconnect_0|rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ;
wire \mm_interconnect_0|spill_enable_s1_agent|m0_write~combout ;
wire \mm_interconnect_0|spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ;
wire \mm_interconnect_0|spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ;
wire \mm_interconnect_0|spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ;
wire \mm_interconnect_0|tick_in_s1_agent|m0_write~combout ;
wire \mm_interconnect_0|tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ;
wire \mm_interconnect_0|tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ;
wire \mm_interconnect_0|tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ;
wire \mm_interconnect_0|time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ;
wire \mm_interconnect_0|time_in_s1_agent|m0_write~combout ;
wire \mm_interconnect_0|time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ;
wire \mm_interconnect_0|time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ;
wire \mm_interconnect_0|time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[1]~q ;
wire \mm_interconnect_0|time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[2]~q ;
wire \mm_interconnect_0|time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[3]~q ;
wire \mm_interconnect_0|time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[4]~q ;
wire \mm_interconnect_0|time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[5]~q ;
wire \mm_interconnect_0|time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[6]~q ;
wire \mm_interconnect_0|time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[7]~q ;
wire \mm_interconnect_0|tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ;
wire \mm_interconnect_0|tx_clk_div_s1_agent|m0_write~combout ;
wire \mm_interconnect_0|tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ;
wire \mm_interconnect_0|tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ;
wire \mm_interconnect_0|tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[1]~q ;
wire \mm_interconnect_0|tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[2]~q ;
wire \mm_interconnect_0|tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[3]~q ;
wire \mm_interconnect_0|tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[4]~q ;
wire \mm_interconnect_0|tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[5]~q ;
wire \mm_interconnect_0|tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[6]~q ;
wire \mm_interconnect_0|wr_data_s1_agent|m0_write~combout ;
wire \mm_interconnect_0|wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ;
wire \mm_interconnect_0|wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ;
wire \mm_interconnect_0|wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ;
wire \rst_controller_001|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \autostart|readdata[0]~0_combout ;
wire \tx_clk_div|readdata[0]~combout ;
wire \currentstate|readdata[0]~q ;
wire \data_o|readdata[0]~q ;
wire \tx_full|readdata[0]~q ;
wire \flags|readdata[0]~q ;
wire \time_out|readdata[0]~q ;
wire \tick_out|readdata[0]~q ;
wire \rx_empty|readdata[0]~q ;
wire \link_start|readdata[0]~0_combout ;
wire \link_disable|readdata[0]~0_combout ;
wire \wr_data|readdata[0]~0_combout ;
wire \rd_data|readdata[0]~0_combout ;
wire \tick_in|readdata[0]~0_combout ;
wire \spill_enable|readdata[0]~0_combout ;
wire \data_i|readdata[0]~combout ;
wire \time_in|readdata[0]~combout ;
wire \currentstate|readdata[1]~q ;
wire \data_i|readdata[1]~combout ;
wire \time_out|readdata[1]~q ;
wire \data_o|readdata[1]~q ;
wire \flags|readdata[1]~q ;
wire \time_in|readdata[1]~combout ;
wire \tx_clk_div|readdata[1]~combout ;
wire \currentstate|readdata[2]~q ;
wire \data_i|readdata[2]~combout ;
wire \time_out|readdata[2]~q ;
wire \data_o|readdata[2]~q ;
wire \flags|readdata[2]~q ;
wire \time_in|readdata[2]~combout ;
wire \tx_clk_div|readdata[2]~combout ;
wire \flags|readdata[3]~q ;
wire \data_i|readdata[3]~combout ;
wire \time_out|readdata[3]~q ;
wire \data_o|readdata[3]~q ;
wire \time_in|readdata[3]~combout ;
wire \tx_clk_div|readdata[3]~combout ;
wire \flags|readdata[4]~q ;
wire \data_i|readdata[4]~combout ;
wire \time_out|readdata[4]~q ;
wire \data_o|readdata[4]~q ;
wire \time_in|readdata[4]~combout ;
wire \tx_clk_div|readdata[4]~combout ;
wire \flags|readdata[5]~q ;
wire \data_i|readdata[5]~combout ;
wire \time_out|readdata[5]~q ;
wire \data_o|readdata[5]~q ;
wire \time_in|readdata[5]~combout ;
wire \tx_clk_div|readdata[5]~combout ;
wire \flags|readdata[6]~q ;
wire \data_i|readdata[6]~combout ;
wire \time_out|readdata[6]~q ;
wire \data_o|readdata[6]~q ;
wire \time_in|readdata[6]~combout ;
wire \tx_clk_div|readdata[6]~combout ;
wire \flags|readdata[7]~q ;
wire \data_i|readdata[7]~combout ;
wire \time_in|readdata[7]~combout ;
wire \time_out|readdata[7]~q ;
wire \data_o|readdata[7]~q ;
wire \data_i|readdata[8]~combout ;
wire \flags|readdata[8]~q ;
wire \data_o|readdata[8]~q ;
wire \flags|readdata[9]~q ;
wire \flags|readdata[10]~q ;
wire \mm_interconnect_0|currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ;
wire \mm_interconnect_0|currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ;
wire \mm_interconnect_0|data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ;
wire \mm_interconnect_0|data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ;
wire \mm_interconnect_0|tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ;
wire \mm_interconnect_0|tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ;
wire \mm_interconnect_0|flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ;
wire \mm_interconnect_0|flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ;
wire \mm_interconnect_0|time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ;
wire \mm_interconnect_0|time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ;
wire \mm_interconnect_0|tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ;
wire \mm_interconnect_0|tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ;
wire \mm_interconnect_0|rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ;
wire \mm_interconnect_0|rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ;
wire \clk_clk~input_o ;
wire \reset_reset_n~input_o ;
wire \currentstate_external_connection_export[0]~input_o ;
wire \data_o_external_connection_export[0]~input_o ;
wire \tx_full_external_connection_export~input_o ;
wire \flags_external_connection_export[0]~input_o ;
wire \time_out_external_connection_export[0]~input_o ;
wire \tick_out_external_connection_export~input_o ;
wire \rx_empty_external_connection_export~input_o ;
wire \currentstate_external_connection_export[1]~input_o ;
wire \time_out_external_connection_export[1]~input_o ;
wire \data_o_external_connection_export[1]~input_o ;
wire \flags_external_connection_export[1]~input_o ;
wire \currentstate_external_connection_export[2]~input_o ;
wire \time_out_external_connection_export[2]~input_o ;
wire \data_o_external_connection_export[2]~input_o ;
wire \flags_external_connection_export[2]~input_o ;
wire \flags_external_connection_export[3]~input_o ;
wire \time_out_external_connection_export[3]~input_o ;
wire \data_o_external_connection_export[3]~input_o ;
wire \flags_external_connection_export[4]~input_o ;
wire \time_out_external_connection_export[4]~input_o ;
wire \data_o_external_connection_export[4]~input_o ;
wire \flags_external_connection_export[5]~input_o ;
wire \time_out_external_connection_export[5]~input_o ;
wire \data_o_external_connection_export[5]~input_o ;
wire \flags_external_connection_export[6]~input_o ;
wire \time_out_external_connection_export[6]~input_o ;
wire \data_o_external_connection_export[6]~input_o ;
wire \flags_external_connection_export[7]~input_o ;
wire \time_out_external_connection_export[7]~input_o ;
wire \data_o_external_connection_export[7]~input_o ;
wire \flags_external_connection_export[8]~input_o ;
wire \data_o_external_connection_export[8]~input_o ;
wire \flags_external_connection_export[9]~input_o ;
wire \flags_external_connection_export[10]~input_o ;


spw_babasu_altera_reset_controller_1 rst_controller_001(
	.h2f_rst_n_0(\hps_0|fpga_interfaces|h2f_rst_n[0] ),
	.altera_reset_synchronizer_int_chain_out(\rst_controller_001|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.clk_clk(\clk_clk~input_o ));

spw_babasu_altera_reset_controller rst_controller(
	.altera_reset_synchronizer_int_chain_out(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.clk_clk(\clk_clk~input_o ),
	.reset_reset_n(\reset_reset_n~input_o ));

spw_babasu_spw_babasu_RX_EMPTY rx_empty(
	.altera_reset_synchronizer_int_chain_out(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.readdata_0(\rx_empty|readdata[0]~q ),
	.int_nxt_addr_reg_dly_3(\mm_interconnect_0|rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_2(\mm_interconnect_0|rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.clk_clk(\clk_clk~input_o ),
	.rx_empty_external_connection_export(\rx_empty_external_connection_export~input_o ));

spw_babasu_spw_babasu_AUTOSTART_3 rd_data(
	.data_out1(\rd_data|data_out~q ),
	.wait_latency_counter_1(\mm_interconnect_0|rd_data_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\mm_interconnect_0|rd_data_s1_translator|wait_latency_counter[0]~q ),
	.reset_n(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.m0_write(\mm_interconnect_0|rd_data_s1_agent|m0_write~combout ),
	.in_data_reg_0(\mm_interconnect_0|rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ),
	.int_nxt_addr_reg_dly_3(\mm_interconnect_0|rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_2(\mm_interconnect_0|rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.readdata_0(\rd_data|readdata[0]~0_combout ),
	.clk(\clk_clk~input_o ));

spw_babasu_spw_babasu_AUTOSTART_2 link_start(
	.data_out1(\link_start|data_out~q ),
	.wait_latency_counter_1(\mm_interconnect_0|link_start_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\mm_interconnect_0|link_start_s1_translator|wait_latency_counter[0]~q ),
	.reset_n(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.m0_write(\mm_interconnect_0|link_start_s1_agent|m0_write~combout ),
	.in_data_reg_0(\mm_interconnect_0|link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ),
	.int_nxt_addr_reg_dly_3(\mm_interconnect_0|link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_2(\mm_interconnect_0|link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.readdata_0(\link_start|readdata[0]~0_combout ),
	.clk(\clk_clk~input_o ));

spw_babasu_spw_babasu_AUTOSTART_1 link_disable(
	.data_out1(\link_disable|data_out~q ),
	.wait_latency_counter_1(\mm_interconnect_0|link_disable_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\mm_interconnect_0|link_disable_s1_translator|wait_latency_counter[0]~q ),
	.reset_n(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.m0_write(\mm_interconnect_0|link_disable_s1_agent|m0_write~combout ),
	.in_data_reg_0(\mm_interconnect_0|link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ),
	.int_nxt_addr_reg_dly_3(\mm_interconnect_0|link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_2(\mm_interconnect_0|link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.readdata_0(\link_disable|readdata[0]~0_combout ),
	.clk(\clk_clk~input_o ));

spw_babasu_spw_babasu_FLAGS flags(
	.altera_reset_synchronizer_int_chain_out(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.readdata_0(\flags|readdata[0]~q ),
	.readdata_1(\flags|readdata[1]~q ),
	.readdata_2(\flags|readdata[2]~q ),
	.readdata_3(\flags|readdata[3]~q ),
	.readdata_4(\flags|readdata[4]~q ),
	.readdata_5(\flags|readdata[5]~q ),
	.readdata_6(\flags|readdata[6]~q ),
	.readdata_7(\flags|readdata[7]~q ),
	.readdata_8(\flags|readdata[8]~q ),
	.readdata_9(\flags|readdata[9]~q ),
	.readdata_10(\flags|readdata[10]~q ),
	.int_nxt_addr_reg_dly_3(\mm_interconnect_0|flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_2(\mm_interconnect_0|flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.clk_clk(\clk_clk~input_o ),
	.flags_external_connection_export_0(\flags_external_connection_export[0]~input_o ),
	.flags_external_connection_export_1(\flags_external_connection_export[1]~input_o ),
	.flags_external_connection_export_2(\flags_external_connection_export[2]~input_o ),
	.flags_external_connection_export_3(\flags_external_connection_export[3]~input_o ),
	.flags_external_connection_export_4(\flags_external_connection_export[4]~input_o ),
	.flags_external_connection_export_5(\flags_external_connection_export[5]~input_o ),
	.flags_external_connection_export_6(\flags_external_connection_export[6]~input_o ),
	.flags_external_connection_export_7(\flags_external_connection_export[7]~input_o ),
	.flags_external_connection_export_8(\flags_external_connection_export[8]~input_o ),
	.flags_external_connection_export_9(\flags_external_connection_export[9]~input_o ),
	.flags_external_connection_export_10(\flags_external_connection_export[10]~input_o ));

spw_babasu_spw_babasu_DATA_O data_o(
	.altera_reset_synchronizer_int_chain_out(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.readdata_0(\data_o|readdata[0]~q ),
	.readdata_1(\data_o|readdata[1]~q ),
	.readdata_2(\data_o|readdata[2]~q ),
	.readdata_3(\data_o|readdata[3]~q ),
	.readdata_4(\data_o|readdata[4]~q ),
	.readdata_5(\data_o|readdata[5]~q ),
	.readdata_6(\data_o|readdata[6]~q ),
	.readdata_7(\data_o|readdata[7]~q ),
	.readdata_8(\data_o|readdata[8]~q ),
	.int_nxt_addr_reg_dly_3(\mm_interconnect_0|data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_2(\mm_interconnect_0|data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.clk_clk(\clk_clk~input_o ),
	.data_o_external_connection_export_0(\data_o_external_connection_export[0]~input_o ),
	.data_o_external_connection_export_1(\data_o_external_connection_export[1]~input_o ),
	.data_o_external_connection_export_2(\data_o_external_connection_export[2]~input_o ),
	.data_o_external_connection_export_3(\data_o_external_connection_export[3]~input_o ),
	.data_o_external_connection_export_4(\data_o_external_connection_export[4]~input_o ),
	.data_o_external_connection_export_5(\data_o_external_connection_export[5]~input_o ),
	.data_o_external_connection_export_6(\data_o_external_connection_export[6]~input_o ),
	.data_o_external_connection_export_7(\data_o_external_connection_export[7]~input_o ),
	.data_o_external_connection_export_8(\data_o_external_connection_export[8]~input_o ));

spw_babasu_spw_babasu_DATA_I data_i(
	.data_out_0(\data_i|data_out[0]~q ),
	.data_out_1(\data_i|data_out[1]~q ),
	.data_out_2(\data_i|data_out[2]~q ),
	.data_out_3(\data_i|data_out[3]~q ),
	.data_out_4(\data_i|data_out[4]~q ),
	.data_out_5(\data_i|data_out[5]~q ),
	.data_out_6(\data_i|data_out[6]~q ),
	.data_out_7(\data_i|data_out[7]~q ),
	.data_out_8(\data_i|data_out[8]~q ),
	.wait_latency_counter_1(\mm_interconnect_0|data_i_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\mm_interconnect_0|data_i_s1_translator|wait_latency_counter[0]~q ),
	.reset_n(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.writedata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mm_interconnect_0|data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[8]~q ,
\mm_interconnect_0|data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[7]~q ,\mm_interconnect_0|data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[6]~q ,
\mm_interconnect_0|data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[5]~q ,\mm_interconnect_0|data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[4]~q ,
\mm_interconnect_0|data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[3]~q ,\mm_interconnect_0|data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[2]~q ,
\mm_interconnect_0|data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[1]~q ,\mm_interconnect_0|data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q }),
	.m0_write(\mm_interconnect_0|data_i_s1_agent|m0_write~combout ),
	.int_nxt_addr_reg_dly_3(\mm_interconnect_0|data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_2(\mm_interconnect_0|data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.readdata_0(\data_i|readdata[0]~combout ),
	.readdata_1(\data_i|readdata[1]~combout ),
	.readdata_2(\data_i|readdata[2]~combout ),
	.readdata_3(\data_i|readdata[3]~combout ),
	.readdata_4(\data_i|readdata[4]~combout ),
	.readdata_5(\data_i|readdata[5]~combout ),
	.readdata_6(\data_i|readdata[6]~combout ),
	.readdata_7(\data_i|readdata[7]~combout ),
	.readdata_8(\data_i|readdata[8]~combout ),
	.clk(\clk_clk~input_o ));

spw_babasu_spw_babasu_CURRENTSTATE currentstate(
	.altera_reset_synchronizer_int_chain_out(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.readdata_0(\currentstate|readdata[0]~q ),
	.readdata_1(\currentstate|readdata[1]~q ),
	.readdata_2(\currentstate|readdata[2]~q ),
	.int_nxt_addr_reg_dly_3(\mm_interconnect_0|currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_2(\mm_interconnect_0|currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.clk_clk(\clk_clk~input_o ),
	.currentstate_external_connection_export_0(\currentstate_external_connection_export[0]~input_o ),
	.currentstate_external_connection_export_1(\currentstate_external_connection_export[1]~input_o ),
	.currentstate_external_connection_export_2(\currentstate_external_connection_export[2]~input_o ));

spw_babasu_spw_babasu_AUTOSTART autostart(
	.data_out1(\autostart|data_out~q ),
	.wait_latency_counter_1(\mm_interconnect_0|autostart_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\mm_interconnect_0|autostart_s1_translator|wait_latency_counter[0]~q ),
	.m0_write(\mm_interconnect_0|autostart_s1_agent|m0_write~combout ),
	.in_data_reg_0(\mm_interconnect_0|autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ),
	.int_nxt_addr_reg_dly_3(\mm_interconnect_0|autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_2(\mm_interconnect_0|autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.reset_n(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.readdata_0(\autostart|readdata[0]~0_combout ),
	.clk(\clk_clk~input_o ));

spw_babasu_spw_babasu_hps_0 hps_0(
	.h2f_rst_n_0(\hps_0|fpga_interfaces|h2f_rst_n[0] ),
	.h2f_ARVALID_0(\hps_0|fpga_interfaces|h2f_ARVALID[0] ),
	.h2f_AWVALID_0(\hps_0|fpga_interfaces|h2f_AWVALID[0] ),
	.h2f_BREADY_0(\hps_0|fpga_interfaces|h2f_BREADY[0] ),
	.h2f_RREADY_0(\hps_0|fpga_interfaces|h2f_RREADY[0] ),
	.h2f_WLAST_0(\hps_0|fpga_interfaces|h2f_WLAST[0] ),
	.h2f_WVALID_0(\hps_0|fpga_interfaces|h2f_WVALID[0] ),
	.h2f_ARADDR_0(\hps_0|fpga_interfaces|h2f_ARADDR[0] ),
	.h2f_ARADDR_1(\hps_0|fpga_interfaces|h2f_ARADDR[1] ),
	.h2f_ARADDR_2(\hps_0|fpga_interfaces|h2f_ARADDR[2] ),
	.h2f_ARADDR_3(\hps_0|fpga_interfaces|h2f_ARADDR[3] ),
	.h2f_ARADDR_4(\hps_0|fpga_interfaces|h2f_ARADDR[4] ),
	.h2f_ARADDR_5(\hps_0|fpga_interfaces|h2f_ARADDR[5] ),
	.h2f_ARADDR_6(\hps_0|fpga_interfaces|h2f_ARADDR[6] ),
	.h2f_ARADDR_7(\hps_0|fpga_interfaces|h2f_ARADDR[7] ),
	.h2f_ARADDR_8(\hps_0|fpga_interfaces|h2f_ARADDR[8] ),
	.h2f_ARBURST_0(\hps_0|fpga_interfaces|h2f_ARBURST[0] ),
	.h2f_ARBURST_1(\hps_0|fpga_interfaces|h2f_ARBURST[1] ),
	.h2f_ARID_0(\hps_0|fpga_interfaces|h2f_ARID[0] ),
	.h2f_ARID_1(\hps_0|fpga_interfaces|h2f_ARID[1] ),
	.h2f_ARID_2(\hps_0|fpga_interfaces|h2f_ARID[2] ),
	.h2f_ARID_3(\hps_0|fpga_interfaces|h2f_ARID[3] ),
	.h2f_ARID_4(\hps_0|fpga_interfaces|h2f_ARID[4] ),
	.h2f_ARID_5(\hps_0|fpga_interfaces|h2f_ARID[5] ),
	.h2f_ARID_6(\hps_0|fpga_interfaces|h2f_ARID[6] ),
	.h2f_ARID_7(\hps_0|fpga_interfaces|h2f_ARID[7] ),
	.h2f_ARID_8(\hps_0|fpga_interfaces|h2f_ARID[8] ),
	.h2f_ARID_9(\hps_0|fpga_interfaces|h2f_ARID[9] ),
	.h2f_ARID_10(\hps_0|fpga_interfaces|h2f_ARID[10] ),
	.h2f_ARID_11(\hps_0|fpga_interfaces|h2f_ARID[11] ),
	.h2f_ARLEN_0(\hps_0|fpga_interfaces|h2f_ARLEN[0] ),
	.h2f_ARLEN_1(\hps_0|fpga_interfaces|h2f_ARLEN[1] ),
	.h2f_ARLEN_2(\hps_0|fpga_interfaces|h2f_ARLEN[2] ),
	.h2f_ARLEN_3(\hps_0|fpga_interfaces|h2f_ARLEN[3] ),
	.h2f_ARSIZE_0(\hps_0|fpga_interfaces|h2f_ARSIZE[0] ),
	.h2f_ARSIZE_1(\hps_0|fpga_interfaces|h2f_ARSIZE[1] ),
	.h2f_ARSIZE_2(\hps_0|fpga_interfaces|h2f_ARSIZE[2] ),
	.h2f_AWADDR_0(\hps_0|fpga_interfaces|h2f_AWADDR[0] ),
	.h2f_AWADDR_1(\hps_0|fpga_interfaces|h2f_AWADDR[1] ),
	.h2f_AWADDR_2(\hps_0|fpga_interfaces|h2f_AWADDR[2] ),
	.h2f_AWADDR_3(\hps_0|fpga_interfaces|h2f_AWADDR[3] ),
	.h2f_AWADDR_4(\hps_0|fpga_interfaces|h2f_AWADDR[4] ),
	.h2f_AWADDR_5(\hps_0|fpga_interfaces|h2f_AWADDR[5] ),
	.h2f_AWADDR_6(\hps_0|fpga_interfaces|h2f_AWADDR[6] ),
	.h2f_AWADDR_7(\hps_0|fpga_interfaces|h2f_AWADDR[7] ),
	.h2f_AWADDR_8(\hps_0|fpga_interfaces|h2f_AWADDR[8] ),
	.h2f_AWBURST_0(\hps_0|fpga_interfaces|h2f_AWBURST[0] ),
	.h2f_AWBURST_1(\hps_0|fpga_interfaces|h2f_AWBURST[1] ),
	.h2f_AWID_0(\hps_0|fpga_interfaces|h2f_AWID[0] ),
	.h2f_AWID_1(\hps_0|fpga_interfaces|h2f_AWID[1] ),
	.h2f_AWID_2(\hps_0|fpga_interfaces|h2f_AWID[2] ),
	.h2f_AWID_3(\hps_0|fpga_interfaces|h2f_AWID[3] ),
	.h2f_AWID_4(\hps_0|fpga_interfaces|h2f_AWID[4] ),
	.h2f_AWID_5(\hps_0|fpga_interfaces|h2f_AWID[5] ),
	.h2f_AWID_6(\hps_0|fpga_interfaces|h2f_AWID[6] ),
	.h2f_AWID_7(\hps_0|fpga_interfaces|h2f_AWID[7] ),
	.h2f_AWID_8(\hps_0|fpga_interfaces|h2f_AWID[8] ),
	.h2f_AWID_9(\hps_0|fpga_interfaces|h2f_AWID[9] ),
	.h2f_AWID_10(\hps_0|fpga_interfaces|h2f_AWID[10] ),
	.h2f_AWID_11(\hps_0|fpga_interfaces|h2f_AWID[11] ),
	.h2f_AWLEN_0(\hps_0|fpga_interfaces|h2f_AWLEN[0] ),
	.h2f_AWLEN_1(\hps_0|fpga_interfaces|h2f_AWLEN[1] ),
	.h2f_AWLEN_2(\hps_0|fpga_interfaces|h2f_AWLEN[2] ),
	.h2f_AWLEN_3(\hps_0|fpga_interfaces|h2f_AWLEN[3] ),
	.h2f_AWSIZE_0(\hps_0|fpga_interfaces|h2f_AWSIZE[0] ),
	.h2f_AWSIZE_1(\hps_0|fpga_interfaces|h2f_AWSIZE[1] ),
	.h2f_AWSIZE_2(\hps_0|fpga_interfaces|h2f_AWSIZE[2] ),
	.h2f_WDATA_0(\hps_0|fpga_interfaces|h2f_WDATA[0] ),
	.h2f_WDATA_1(\hps_0|fpga_interfaces|h2f_WDATA[1] ),
	.h2f_WDATA_2(\hps_0|fpga_interfaces|h2f_WDATA[2] ),
	.h2f_WDATA_3(\hps_0|fpga_interfaces|h2f_WDATA[3] ),
	.h2f_WDATA_4(\hps_0|fpga_interfaces|h2f_WDATA[4] ),
	.h2f_WDATA_5(\hps_0|fpga_interfaces|h2f_WDATA[5] ),
	.h2f_WDATA_6(\hps_0|fpga_interfaces|h2f_WDATA[6] ),
	.h2f_WDATA_7(\hps_0|fpga_interfaces|h2f_WDATA[7] ),
	.h2f_WDATA_8(\hps_0|fpga_interfaces|h2f_WDATA[8] ),
	.h2f_WSTRB_0(\hps_0|fpga_interfaces|h2f_WSTRB[0] ),
	.h2f_WSTRB_1(\hps_0|fpga_interfaces|h2f_WSTRB[1] ),
	.h2f_WSTRB_2(\hps_0|fpga_interfaces|h2f_WSTRB[2] ),
	.h2f_WSTRB_3(\hps_0|fpga_interfaces|h2f_WSTRB[3] ),
	.cmd_sink_ready(\mm_interconnect_0|hps_0_h2f_axi_master_rd_limiter|cmd_sink_ready~0_combout ),
	.nonposted_cmd_accepted(\mm_interconnect_0|hps_0_h2f_axi_master_wr_limiter|nonposted_cmd_accepted~0_combout ),
	.WideOr1(\mm_interconnect_0|rsp_mux|WideOr1~combout ),
	.src_payload_0(\mm_interconnect_0|rsp_mux_001|src_payload[0]~combout ),
	.WideOr11(\mm_interconnect_0|rsp_mux_001|WideOr1~combout ),
	.nonposted_cmd_accepted1(\mm_interconnect_0|hps_0_h2f_axi_master_wr_limiter|nonposted_cmd_accepted~1_combout ),
	.src_data_105(\mm_interconnect_0|rsp_mux|src_data[105]~combout ),
	.src_data_106(\mm_interconnect_0|rsp_mux|src_data[106]~combout ),
	.src_data_107(\mm_interconnect_0|rsp_mux|src_data[107]~combout ),
	.src_data_108(\mm_interconnect_0|rsp_mux|src_data[108]~combout ),
	.src_data_109(\mm_interconnect_0|rsp_mux|src_data[109]~combout ),
	.src_data_110(\mm_interconnect_0|rsp_mux|src_data[110]~combout ),
	.src_data_111(\mm_interconnect_0|rsp_mux|src_data[111]~combout ),
	.src_data_112(\mm_interconnect_0|rsp_mux|src_data[112]~combout ),
	.src_data_113(\mm_interconnect_0|rsp_mux|src_data[113]~combout ),
	.src_data_114(\mm_interconnect_0|rsp_mux|src_data[114]~combout ),
	.src_data_115(\mm_interconnect_0|rsp_mux|src_data[115]~combout ),
	.src_data_116(\mm_interconnect_0|rsp_mux|src_data[116]~combout ),
	.src_data_0(\mm_interconnect_0|rsp_mux_001|src_data[0]~20_combout ),
	.src_payload(\mm_interconnect_0|rsp_mux_001|src_payload~30_combout ),
	.src_payload1(\mm_interconnect_0|rsp_mux_001|src_payload~38_combout ),
	.src_payload2(\mm_interconnect_0|rsp_mux_001|src_payload~45_combout ),
	.src_payload3(\mm_interconnect_0|rsp_mux_001|src_payload~52_combout ),
	.src_payload4(\mm_interconnect_0|rsp_mux_001|src_payload~59_combout ),
	.src_payload5(\mm_interconnect_0|rsp_mux_001|src_payload~66_combout ),
	.src_payload6(\mm_interconnect_0|rsp_mux_001|src_payload~72_combout ),
	.src_payload7(\mm_interconnect_0|rsp_mux_001|src_payload~75_combout ),
	.src_payload8(\mm_interconnect_0|rsp_mux_001|src_payload~76_combout ),
	.src_payload9(\mm_interconnect_0|rsp_mux_001|src_payload~77_combout ),
	.src_data_1051(\mm_interconnect_0|rsp_mux_001|src_data[105]~combout ),
	.src_data_1061(\mm_interconnect_0|rsp_mux_001|src_data[106]~combout ),
	.src_data_1071(\mm_interconnect_0|rsp_mux_001|src_data[107]~combout ),
	.src_data_1081(\mm_interconnect_0|rsp_mux_001|src_data[108]~combout ),
	.src_data_1091(\mm_interconnect_0|rsp_mux_001|src_data[109]~combout ),
	.src_data_1101(\mm_interconnect_0|rsp_mux_001|src_data[110]~combout ),
	.src_data_1111(\mm_interconnect_0|rsp_mux_001|src_data[111]~combout ),
	.src_data_1121(\mm_interconnect_0|rsp_mux_001|src_data[112]~combout ),
	.src_data_1131(\mm_interconnect_0|rsp_mux_001|src_data[113]~combout ),
	.src_data_1141(\mm_interconnect_0|rsp_mux_001|src_data[114]~combout ),
	.src_data_1151(\mm_interconnect_0|rsp_mux_001|src_data[115]~combout ),
	.src_data_1161(\mm_interconnect_0|rsp_mux_001|src_data[116]~combout ),
	.clk_clk(\clk_clk~input_o ));

spw_babasu_spw_babasu_AUTOSTART_6 wr_data(
	.data_out1(\wr_data|data_out~q ),
	.wait_latency_counter_1(\mm_interconnect_0|wr_data_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\mm_interconnect_0|wr_data_s1_translator|wait_latency_counter[0]~q ),
	.reset_n(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.m0_write(\mm_interconnect_0|wr_data_s1_agent|m0_write~combout ),
	.in_data_reg_0(\mm_interconnect_0|wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ),
	.int_nxt_addr_reg_dly_3(\mm_interconnect_0|wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_2(\mm_interconnect_0|wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.readdata_0(\wr_data|readdata[0]~0_combout ),
	.clk(\clk_clk~input_o ));

spw_babasu_spw_babasu_RX_EMPTY_2 tx_full(
	.altera_reset_synchronizer_int_chain_out(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.readdata_0(\tx_full|readdata[0]~q ),
	.int_nxt_addr_reg_dly_3(\mm_interconnect_0|tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_2(\mm_interconnect_0|tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.clk_clk(\clk_clk~input_o ),
	.tx_full_external_connection_export(\tx_full_external_connection_export~input_o ));

spw_babasu_spw_babasu_TX_CLK_DIV tx_clk_div(
	.data_out_0(\tx_clk_div|data_out[0]~q ),
	.data_out_1(\tx_clk_div|data_out[1]~q ),
	.data_out_2(\tx_clk_div|data_out[2]~q ),
	.data_out_3(\tx_clk_div|data_out[3]~q ),
	.data_out_4(\tx_clk_div|data_out[4]~q ),
	.data_out_5(\tx_clk_div|data_out[5]~q ),
	.data_out_6(\tx_clk_div|data_out[6]~q ),
	.wait_latency_counter_1(\mm_interconnect_0|tx_clk_div_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\mm_interconnect_0|tx_clk_div_s1_translator|wait_latency_counter[0]~q ),
	.reset_n(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.in_data_reg_0(\mm_interconnect_0|tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ),
	.m0_write(\mm_interconnect_0|tx_clk_div_s1_agent|m0_write~combout ),
	.int_nxt_addr_reg_dly_3(\mm_interconnect_0|tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_2(\mm_interconnect_0|tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.in_data_reg_1(\mm_interconnect_0|tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[1]~q ),
	.writedata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mm_interconnect_0|tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[6]~q ,
\mm_interconnect_0|tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[5]~q ,\mm_interconnect_0|tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[4]~q ,
\mm_interconnect_0|tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[3]~q ,\mm_interconnect_0|tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[2]~q ,gnd,gnd}),
	.readdata_0(\tx_clk_div|readdata[0]~combout ),
	.readdata_1(\tx_clk_div|readdata[1]~combout ),
	.readdata_2(\tx_clk_div|readdata[2]~combout ),
	.readdata_3(\tx_clk_div|readdata[3]~combout ),
	.readdata_4(\tx_clk_div|readdata[4]~combout ),
	.readdata_5(\tx_clk_div|readdata[5]~combout ),
	.readdata_6(\tx_clk_div|readdata[6]~combout ),
	.clk(\clk_clk~input_o ));

spw_babasu_spw_babasu_TIME_OUT time_out(
	.altera_reset_synchronizer_int_chain_out(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.readdata_0(\time_out|readdata[0]~q ),
	.readdata_1(\time_out|readdata[1]~q ),
	.readdata_2(\time_out|readdata[2]~q ),
	.readdata_3(\time_out|readdata[3]~q ),
	.readdata_4(\time_out|readdata[4]~q ),
	.readdata_5(\time_out|readdata[5]~q ),
	.readdata_6(\time_out|readdata[6]~q ),
	.readdata_7(\time_out|readdata[7]~q ),
	.int_nxt_addr_reg_dly_3(\mm_interconnect_0|time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_2(\mm_interconnect_0|time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.clk_clk(\clk_clk~input_o ),
	.time_out_external_connection_export_0(\time_out_external_connection_export[0]~input_o ),
	.time_out_external_connection_export_1(\time_out_external_connection_export[1]~input_o ),
	.time_out_external_connection_export_2(\time_out_external_connection_export[2]~input_o ),
	.time_out_external_connection_export_3(\time_out_external_connection_export[3]~input_o ),
	.time_out_external_connection_export_4(\time_out_external_connection_export[4]~input_o ),
	.time_out_external_connection_export_5(\time_out_external_connection_export[5]~input_o ),
	.time_out_external_connection_export_6(\time_out_external_connection_export[6]~input_o ),
	.time_out_external_connection_export_7(\time_out_external_connection_export[7]~input_o ));

spw_babasu_spw_babasu_TIME_IN time_in(
	.data_out_0(\time_in|data_out[0]~q ),
	.data_out_1(\time_in|data_out[1]~q ),
	.data_out_2(\time_in|data_out[2]~q ),
	.data_out_3(\time_in|data_out[3]~q ),
	.data_out_4(\time_in|data_out[4]~q ),
	.data_out_5(\time_in|data_out[5]~q ),
	.data_out_6(\time_in|data_out[6]~q ),
	.data_out_7(\time_in|data_out[7]~q ),
	.wait_latency_counter_1(\mm_interconnect_0|time_in_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\mm_interconnect_0|time_in_s1_translator|wait_latency_counter[0]~q ),
	.reset_n(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.writedata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mm_interconnect_0|time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[7]~q ,
\mm_interconnect_0|time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[6]~q ,\mm_interconnect_0|time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[5]~q ,
\mm_interconnect_0|time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[4]~q ,\mm_interconnect_0|time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[3]~q ,
\mm_interconnect_0|time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[2]~q ,\mm_interconnect_0|time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[1]~q ,
\mm_interconnect_0|time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q }),
	.m0_write(\mm_interconnect_0|time_in_s1_agent|m0_write~combout ),
	.int_nxt_addr_reg_dly_3(\mm_interconnect_0|time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_2(\mm_interconnect_0|time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.readdata_0(\time_in|readdata[0]~combout ),
	.readdata_1(\time_in|readdata[1]~combout ),
	.readdata_2(\time_in|readdata[2]~combout ),
	.readdata_3(\time_in|readdata[3]~combout ),
	.readdata_4(\time_in|readdata[4]~combout ),
	.readdata_5(\time_in|readdata[5]~combout ),
	.readdata_6(\time_in|readdata[6]~combout ),
	.readdata_7(\time_in|readdata[7]~combout ),
	.clk(\clk_clk~input_o ));

spw_babasu_spw_babasu_RX_EMPTY_1 tick_out(
	.altera_reset_synchronizer_int_chain_out(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.readdata_0(\tick_out|readdata[0]~q ),
	.int_nxt_addr_reg_dly_3(\mm_interconnect_0|tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_2(\mm_interconnect_0|tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.clk_clk(\clk_clk~input_o ),
	.tick_out_external_connection_export(\tick_out_external_connection_export~input_o ));

spw_babasu_spw_babasu_AUTOSTART_5 tick_in(
	.data_out1(\tick_in|data_out~q ),
	.wait_latency_counter_1(\mm_interconnect_0|tick_in_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\mm_interconnect_0|tick_in_s1_translator|wait_latency_counter[0]~q ),
	.reset_n(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.m0_write(\mm_interconnect_0|tick_in_s1_agent|m0_write~combout ),
	.in_data_reg_0(\mm_interconnect_0|tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ),
	.int_nxt_addr_reg_dly_3(\mm_interconnect_0|tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_2(\mm_interconnect_0|tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.readdata_0(\tick_in|readdata[0]~0_combout ),
	.clk(\clk_clk~input_o ));

spw_babasu_spw_babasu_AUTOSTART_4 spill_enable(
	.data_out1(\spill_enable|data_out~q ),
	.wait_latency_counter_1(\mm_interconnect_0|spill_enable_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\mm_interconnect_0|spill_enable_s1_translator|wait_latency_counter[0]~q ),
	.reset_n(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.m0_write(\mm_interconnect_0|spill_enable_s1_agent|m0_write~combout ),
	.in_data_reg_0(\mm_interconnect_0|spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ),
	.int_nxt_addr_reg_dly_3(\mm_interconnect_0|spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_2(\mm_interconnect_0|spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.readdata_0(\spill_enable|readdata[0]~0_combout ),
	.clk(\clk_clk~input_o ));

spw_babasu_spw_babasu_mm_interconnect_0 mm_interconnect_0(
	.h2f_ARVALID_0(\hps_0|fpga_interfaces|h2f_ARVALID[0] ),
	.h2f_AWVALID_0(\hps_0|fpga_interfaces|h2f_AWVALID[0] ),
	.h2f_BREADY_0(\hps_0|fpga_interfaces|h2f_BREADY[0] ),
	.h2f_RREADY_0(\hps_0|fpga_interfaces|h2f_RREADY[0] ),
	.h2f_WLAST_0(\hps_0|fpga_interfaces|h2f_WLAST[0] ),
	.h2f_WVALID_0(\hps_0|fpga_interfaces|h2f_WVALID[0] ),
	.h2f_ARADDR_0(\hps_0|fpga_interfaces|h2f_ARADDR[0] ),
	.h2f_ARADDR_1(\hps_0|fpga_interfaces|h2f_ARADDR[1] ),
	.h2f_ARADDR_2(\hps_0|fpga_interfaces|h2f_ARADDR[2] ),
	.h2f_ARADDR_3(\hps_0|fpga_interfaces|h2f_ARADDR[3] ),
	.h2f_ARADDR_4(\hps_0|fpga_interfaces|h2f_ARADDR[4] ),
	.h2f_ARADDR_5(\hps_0|fpga_interfaces|h2f_ARADDR[5] ),
	.h2f_ARADDR_6(\hps_0|fpga_interfaces|h2f_ARADDR[6] ),
	.h2f_ARADDR_7(\hps_0|fpga_interfaces|h2f_ARADDR[7] ),
	.h2f_ARADDR_8(\hps_0|fpga_interfaces|h2f_ARADDR[8] ),
	.h2f_ARBURST_0(\hps_0|fpga_interfaces|h2f_ARBURST[0] ),
	.h2f_ARBURST_1(\hps_0|fpga_interfaces|h2f_ARBURST[1] ),
	.h2f_ARID_0(\hps_0|fpga_interfaces|h2f_ARID[0] ),
	.h2f_ARID_1(\hps_0|fpga_interfaces|h2f_ARID[1] ),
	.h2f_ARID_2(\hps_0|fpga_interfaces|h2f_ARID[2] ),
	.h2f_ARID_3(\hps_0|fpga_interfaces|h2f_ARID[3] ),
	.h2f_ARID_4(\hps_0|fpga_interfaces|h2f_ARID[4] ),
	.h2f_ARID_5(\hps_0|fpga_interfaces|h2f_ARID[5] ),
	.h2f_ARID_6(\hps_0|fpga_interfaces|h2f_ARID[6] ),
	.h2f_ARID_7(\hps_0|fpga_interfaces|h2f_ARID[7] ),
	.h2f_ARID_8(\hps_0|fpga_interfaces|h2f_ARID[8] ),
	.h2f_ARID_9(\hps_0|fpga_interfaces|h2f_ARID[9] ),
	.h2f_ARID_10(\hps_0|fpga_interfaces|h2f_ARID[10] ),
	.h2f_ARID_11(\hps_0|fpga_interfaces|h2f_ARID[11] ),
	.h2f_ARLEN_0(\hps_0|fpga_interfaces|h2f_ARLEN[0] ),
	.h2f_ARLEN_1(\hps_0|fpga_interfaces|h2f_ARLEN[1] ),
	.h2f_ARLEN_2(\hps_0|fpga_interfaces|h2f_ARLEN[2] ),
	.h2f_ARLEN_3(\hps_0|fpga_interfaces|h2f_ARLEN[3] ),
	.h2f_ARSIZE_0(\hps_0|fpga_interfaces|h2f_ARSIZE[0] ),
	.h2f_ARSIZE_1(\hps_0|fpga_interfaces|h2f_ARSIZE[1] ),
	.h2f_ARSIZE_2(\hps_0|fpga_interfaces|h2f_ARSIZE[2] ),
	.h2f_AWADDR_0(\hps_0|fpga_interfaces|h2f_AWADDR[0] ),
	.h2f_AWADDR_1(\hps_0|fpga_interfaces|h2f_AWADDR[1] ),
	.h2f_AWADDR_2(\hps_0|fpga_interfaces|h2f_AWADDR[2] ),
	.h2f_AWADDR_3(\hps_0|fpga_interfaces|h2f_AWADDR[3] ),
	.h2f_AWADDR_4(\hps_0|fpga_interfaces|h2f_AWADDR[4] ),
	.h2f_AWADDR_5(\hps_0|fpga_interfaces|h2f_AWADDR[5] ),
	.h2f_AWADDR_6(\hps_0|fpga_interfaces|h2f_AWADDR[6] ),
	.h2f_AWADDR_7(\hps_0|fpga_interfaces|h2f_AWADDR[7] ),
	.h2f_AWADDR_8(\hps_0|fpga_interfaces|h2f_AWADDR[8] ),
	.h2f_AWBURST_0(\hps_0|fpga_interfaces|h2f_AWBURST[0] ),
	.h2f_AWBURST_1(\hps_0|fpga_interfaces|h2f_AWBURST[1] ),
	.h2f_AWID_0(\hps_0|fpga_interfaces|h2f_AWID[0] ),
	.h2f_AWID_1(\hps_0|fpga_interfaces|h2f_AWID[1] ),
	.h2f_AWID_2(\hps_0|fpga_interfaces|h2f_AWID[2] ),
	.h2f_AWID_3(\hps_0|fpga_interfaces|h2f_AWID[3] ),
	.h2f_AWID_4(\hps_0|fpga_interfaces|h2f_AWID[4] ),
	.h2f_AWID_5(\hps_0|fpga_interfaces|h2f_AWID[5] ),
	.h2f_AWID_6(\hps_0|fpga_interfaces|h2f_AWID[6] ),
	.h2f_AWID_7(\hps_0|fpga_interfaces|h2f_AWID[7] ),
	.h2f_AWID_8(\hps_0|fpga_interfaces|h2f_AWID[8] ),
	.h2f_AWID_9(\hps_0|fpga_interfaces|h2f_AWID[9] ),
	.h2f_AWID_10(\hps_0|fpga_interfaces|h2f_AWID[10] ),
	.h2f_AWID_11(\hps_0|fpga_interfaces|h2f_AWID[11] ),
	.h2f_AWLEN_0(\hps_0|fpga_interfaces|h2f_AWLEN[0] ),
	.h2f_AWLEN_1(\hps_0|fpga_interfaces|h2f_AWLEN[1] ),
	.h2f_AWLEN_2(\hps_0|fpga_interfaces|h2f_AWLEN[2] ),
	.h2f_AWLEN_3(\hps_0|fpga_interfaces|h2f_AWLEN[3] ),
	.h2f_AWSIZE_0(\hps_0|fpga_interfaces|h2f_AWSIZE[0] ),
	.h2f_AWSIZE_1(\hps_0|fpga_interfaces|h2f_AWSIZE[1] ),
	.h2f_AWSIZE_2(\hps_0|fpga_interfaces|h2f_AWSIZE[2] ),
	.h2f_WDATA_0(\hps_0|fpga_interfaces|h2f_WDATA[0] ),
	.h2f_WDATA_1(\hps_0|fpga_interfaces|h2f_WDATA[1] ),
	.h2f_WDATA_2(\hps_0|fpga_interfaces|h2f_WDATA[2] ),
	.h2f_WDATA_3(\hps_0|fpga_interfaces|h2f_WDATA[3] ),
	.h2f_WDATA_4(\hps_0|fpga_interfaces|h2f_WDATA[4] ),
	.h2f_WDATA_5(\hps_0|fpga_interfaces|h2f_WDATA[5] ),
	.h2f_WDATA_6(\hps_0|fpga_interfaces|h2f_WDATA[6] ),
	.h2f_WDATA_7(\hps_0|fpga_interfaces|h2f_WDATA[7] ),
	.h2f_WDATA_8(\hps_0|fpga_interfaces|h2f_WDATA[8] ),
	.h2f_WSTRB_0(\hps_0|fpga_interfaces|h2f_WSTRB[0] ),
	.h2f_WSTRB_1(\hps_0|fpga_interfaces|h2f_WSTRB[1] ),
	.h2f_WSTRB_2(\hps_0|fpga_interfaces|h2f_WSTRB[2] ),
	.h2f_WSTRB_3(\hps_0|fpga_interfaces|h2f_WSTRB[3] ),
	.wait_latency_counter_1(\mm_interconnect_0|link_disable_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\mm_interconnect_0|link_disable_s1_translator|wait_latency_counter[0]~q ),
	.wait_latency_counter_11(\mm_interconnect_0|tx_clk_div_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_01(\mm_interconnect_0|tx_clk_div_s1_translator|wait_latency_counter[0]~q ),
	.wait_latency_counter_12(\mm_interconnect_0|spill_enable_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_02(\mm_interconnect_0|spill_enable_s1_translator|wait_latency_counter[0]~q ),
	.wait_latency_counter_13(\mm_interconnect_0|tick_in_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_03(\mm_interconnect_0|tick_in_s1_translator|wait_latency_counter[0]~q ),
	.wait_latency_counter_14(\mm_interconnect_0|time_in_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_04(\mm_interconnect_0|time_in_s1_translator|wait_latency_counter[0]~q ),
	.wait_latency_counter_15(\mm_interconnect_0|data_i_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_05(\mm_interconnect_0|data_i_s1_translator|wait_latency_counter[0]~q ),
	.wait_latency_counter_16(\mm_interconnect_0|rd_data_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_06(\mm_interconnect_0|rd_data_s1_translator|wait_latency_counter[0]~q ),
	.wait_latency_counter_17(\mm_interconnect_0|link_start_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_07(\mm_interconnect_0|link_start_s1_translator|wait_latency_counter[0]~q ),
	.wait_latency_counter_18(\mm_interconnect_0|autostart_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_08(\mm_interconnect_0|autostart_s1_translator|wait_latency_counter[0]~q ),
	.wait_latency_counter_19(\mm_interconnect_0|wr_data_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_09(\mm_interconnect_0|wr_data_s1_translator|wait_latency_counter[0]~q ),
	.cmd_sink_ready(\mm_interconnect_0|hps_0_h2f_axi_master_rd_limiter|cmd_sink_ready~0_combout ),
	.nonposted_cmd_accepted(\mm_interconnect_0|hps_0_h2f_axi_master_wr_limiter|nonposted_cmd_accepted~0_combout ),
	.WideOr1(\mm_interconnect_0|rsp_mux|WideOr1~combout ),
	.src_payload_0(\mm_interconnect_0|rsp_mux_001|src_payload[0]~combout ),
	.WideOr11(\mm_interconnect_0|rsp_mux_001|WideOr1~combout ),
	.nonposted_cmd_accepted1(\mm_interconnect_0|hps_0_h2f_axi_master_wr_limiter|nonposted_cmd_accepted~1_combout ),
	.src_data_105(\mm_interconnect_0|rsp_mux|src_data[105]~combout ),
	.src_data_106(\mm_interconnect_0|rsp_mux|src_data[106]~combout ),
	.src_data_107(\mm_interconnect_0|rsp_mux|src_data[107]~combout ),
	.src_data_108(\mm_interconnect_0|rsp_mux|src_data[108]~combout ),
	.src_data_109(\mm_interconnect_0|rsp_mux|src_data[109]~combout ),
	.src_data_110(\mm_interconnect_0|rsp_mux|src_data[110]~combout ),
	.src_data_111(\mm_interconnect_0|rsp_mux|src_data[111]~combout ),
	.src_data_112(\mm_interconnect_0|rsp_mux|src_data[112]~combout ),
	.src_data_113(\mm_interconnect_0|rsp_mux|src_data[113]~combout ),
	.src_data_114(\mm_interconnect_0|rsp_mux|src_data[114]~combout ),
	.src_data_115(\mm_interconnect_0|rsp_mux|src_data[115]~combout ),
	.src_data_116(\mm_interconnect_0|rsp_mux|src_data[116]~combout ),
	.src_data_0(\mm_interconnect_0|rsp_mux_001|src_data[0]~20_combout ),
	.src_payload(\mm_interconnect_0|rsp_mux_001|src_payload~30_combout ),
	.src_payload1(\mm_interconnect_0|rsp_mux_001|src_payload~38_combout ),
	.src_payload2(\mm_interconnect_0|rsp_mux_001|src_payload~45_combout ),
	.src_payload3(\mm_interconnect_0|rsp_mux_001|src_payload~52_combout ),
	.src_payload4(\mm_interconnect_0|rsp_mux_001|src_payload~59_combout ),
	.src_payload5(\mm_interconnect_0|rsp_mux_001|src_payload~66_combout ),
	.src_payload6(\mm_interconnect_0|rsp_mux_001|src_payload~72_combout ),
	.src_payload7(\mm_interconnect_0|rsp_mux_001|src_payload~75_combout ),
	.src_payload8(\mm_interconnect_0|rsp_mux_001|src_payload~76_combout ),
	.src_payload9(\mm_interconnect_0|rsp_mux_001|src_payload~77_combout ),
	.src_data_1051(\mm_interconnect_0|rsp_mux_001|src_data[105]~combout ),
	.src_data_1061(\mm_interconnect_0|rsp_mux_001|src_data[106]~combout ),
	.src_data_1071(\mm_interconnect_0|rsp_mux_001|src_data[107]~combout ),
	.src_data_1081(\mm_interconnect_0|rsp_mux_001|src_data[108]~combout ),
	.src_data_1091(\mm_interconnect_0|rsp_mux_001|src_data[109]~combout ),
	.src_data_1101(\mm_interconnect_0|rsp_mux_001|src_data[110]~combout ),
	.src_data_1111(\mm_interconnect_0|rsp_mux_001|src_data[111]~combout ),
	.src_data_1121(\mm_interconnect_0|rsp_mux_001|src_data[112]~combout ),
	.src_data_1131(\mm_interconnect_0|rsp_mux_001|src_data[113]~combout ),
	.src_data_1141(\mm_interconnect_0|rsp_mux_001|src_data[114]~combout ),
	.src_data_1151(\mm_interconnect_0|rsp_mux_001|src_data[115]~combout ),
	.src_data_1161(\mm_interconnect_0|rsp_mux_001|src_data[116]~combout ),
	.m0_write(\mm_interconnect_0|autostart_s1_agent|m0_write~combout ),
	.in_data_reg_0(\mm_interconnect_0|autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ),
	.int_nxt_addr_reg_dly_3(\mm_interconnect_0|autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_2(\mm_interconnect_0|autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.altera_reset_synchronizer_int_chain_out(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.in_data_reg_01(\mm_interconnect_0|data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ),
	.m0_write1(\mm_interconnect_0|data_i_s1_agent|m0_write~combout ),
	.int_nxt_addr_reg_dly_31(\mm_interconnect_0|data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_21(\mm_interconnect_0|data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.in_data_reg_1(\mm_interconnect_0|data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[1]~q ),
	.in_data_reg_2(\mm_interconnect_0|data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[2]~q ),
	.in_data_reg_3(\mm_interconnect_0|data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[3]~q ),
	.in_data_reg_4(\mm_interconnect_0|data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[4]~q ),
	.in_data_reg_5(\mm_interconnect_0|data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[5]~q ),
	.in_data_reg_6(\mm_interconnect_0|data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[6]~q ),
	.in_data_reg_7(\mm_interconnect_0|data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[7]~q ),
	.in_data_reg_8(\mm_interconnect_0|data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[8]~q ),
	.m0_write2(\mm_interconnect_0|link_disable_s1_agent|m0_write~combout ),
	.in_data_reg_02(\mm_interconnect_0|link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ),
	.int_nxt_addr_reg_dly_32(\mm_interconnect_0|link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_22(\mm_interconnect_0|link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.m0_write3(\mm_interconnect_0|link_start_s1_agent|m0_write~combout ),
	.in_data_reg_03(\mm_interconnect_0|link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ),
	.int_nxt_addr_reg_dly_33(\mm_interconnect_0|link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_23(\mm_interconnect_0|link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.m0_write4(\mm_interconnect_0|rd_data_s1_agent|m0_write~combout ),
	.in_data_reg_04(\mm_interconnect_0|rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ),
	.int_nxt_addr_reg_dly_34(\mm_interconnect_0|rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_24(\mm_interconnect_0|rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.m0_write5(\mm_interconnect_0|spill_enable_s1_agent|m0_write~combout ),
	.in_data_reg_05(\mm_interconnect_0|spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ),
	.int_nxt_addr_reg_dly_35(\mm_interconnect_0|spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_25(\mm_interconnect_0|spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.m0_write6(\mm_interconnect_0|tick_in_s1_agent|m0_write~combout ),
	.in_data_reg_06(\mm_interconnect_0|tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ),
	.int_nxt_addr_reg_dly_36(\mm_interconnect_0|tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_26(\mm_interconnect_0|tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.in_data_reg_07(\mm_interconnect_0|time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ),
	.m0_write7(\mm_interconnect_0|time_in_s1_agent|m0_write~combout ),
	.int_nxt_addr_reg_dly_37(\mm_interconnect_0|time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_27(\mm_interconnect_0|time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.in_data_reg_11(\mm_interconnect_0|time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[1]~q ),
	.in_data_reg_21(\mm_interconnect_0|time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[2]~q ),
	.in_data_reg_31(\mm_interconnect_0|time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[3]~q ),
	.in_data_reg_41(\mm_interconnect_0|time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[4]~q ),
	.in_data_reg_51(\mm_interconnect_0|time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[5]~q ),
	.in_data_reg_61(\mm_interconnect_0|time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[6]~q ),
	.in_data_reg_71(\mm_interconnect_0|time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[7]~q ),
	.in_data_reg_08(\mm_interconnect_0|tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ),
	.m0_write8(\mm_interconnect_0|tx_clk_div_s1_agent|m0_write~combout ),
	.int_nxt_addr_reg_dly_38(\mm_interconnect_0|tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_28(\mm_interconnect_0|tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.in_data_reg_12(\mm_interconnect_0|tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[1]~q ),
	.in_data_reg_22(\mm_interconnect_0|tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[2]~q ),
	.in_data_reg_32(\mm_interconnect_0|tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[3]~q ),
	.in_data_reg_42(\mm_interconnect_0|tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[4]~q ),
	.in_data_reg_52(\mm_interconnect_0|tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[5]~q ),
	.in_data_reg_62(\mm_interconnect_0|tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[6]~q ),
	.m0_write9(\mm_interconnect_0|wr_data_s1_agent|m0_write~combout ),
	.in_data_reg_09(\mm_interconnect_0|wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ),
	.int_nxt_addr_reg_dly_39(\mm_interconnect_0|wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_29(\mm_interconnect_0|wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.altera_reset_synchronizer_int_chain_out1(\rst_controller_001|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.readdata_0(\autostart|readdata[0]~0_combout ),
	.readdata_01(\tx_clk_div|readdata[0]~combout ),
	.readdata_02(\currentstate|readdata[0]~q ),
	.readdata_03(\data_o|readdata[0]~q ),
	.readdata_04(\tx_full|readdata[0]~q ),
	.readdata_05(\flags|readdata[0]~q ),
	.readdata_06(\time_out|readdata[0]~q ),
	.readdata_07(\tick_out|readdata[0]~q ),
	.readdata_08(\rx_empty|readdata[0]~q ),
	.readdata_09(\link_start|readdata[0]~0_combout ),
	.readdata_010(\link_disable|readdata[0]~0_combout ),
	.readdata_011(\wr_data|readdata[0]~0_combout ),
	.readdata_012(\rd_data|readdata[0]~0_combout ),
	.readdata_013(\tick_in|readdata[0]~0_combout ),
	.readdata_014(\spill_enable|readdata[0]~0_combout ),
	.readdata_015(\data_i|readdata[0]~combout ),
	.readdata_016(\time_in|readdata[0]~combout ),
	.readdata_1(\currentstate|readdata[1]~q ),
	.readdata_11(\data_i|readdata[1]~combout ),
	.readdata_12(\time_out|readdata[1]~q ),
	.readdata_13(\data_o|readdata[1]~q ),
	.readdata_14(\flags|readdata[1]~q ),
	.readdata_15(\time_in|readdata[1]~combout ),
	.readdata_16(\tx_clk_div|readdata[1]~combout ),
	.readdata_2(\currentstate|readdata[2]~q ),
	.readdata_21(\data_i|readdata[2]~combout ),
	.readdata_22(\time_out|readdata[2]~q ),
	.readdata_23(\data_o|readdata[2]~q ),
	.readdata_24(\flags|readdata[2]~q ),
	.readdata_25(\time_in|readdata[2]~combout ),
	.readdata_26(\tx_clk_div|readdata[2]~combout ),
	.readdata_3(\flags|readdata[3]~q ),
	.readdata_31(\data_i|readdata[3]~combout ),
	.readdata_32(\time_out|readdata[3]~q ),
	.readdata_33(\data_o|readdata[3]~q ),
	.readdata_34(\time_in|readdata[3]~combout ),
	.readdata_35(\tx_clk_div|readdata[3]~combout ),
	.readdata_4(\flags|readdata[4]~q ),
	.readdata_41(\data_i|readdata[4]~combout ),
	.readdata_42(\time_out|readdata[4]~q ),
	.readdata_43(\data_o|readdata[4]~q ),
	.readdata_44(\time_in|readdata[4]~combout ),
	.readdata_45(\tx_clk_div|readdata[4]~combout ),
	.readdata_5(\flags|readdata[5]~q ),
	.readdata_51(\data_i|readdata[5]~combout ),
	.readdata_52(\time_out|readdata[5]~q ),
	.readdata_53(\data_o|readdata[5]~q ),
	.readdata_54(\time_in|readdata[5]~combout ),
	.readdata_55(\tx_clk_div|readdata[5]~combout ),
	.readdata_6(\flags|readdata[6]~q ),
	.readdata_61(\data_i|readdata[6]~combout ),
	.readdata_62(\time_out|readdata[6]~q ),
	.readdata_63(\data_o|readdata[6]~q ),
	.readdata_64(\time_in|readdata[6]~combout ),
	.readdata_65(\tx_clk_div|readdata[6]~combout ),
	.readdata_7(\flags|readdata[7]~q ),
	.readdata_71(\data_i|readdata[7]~combout ),
	.readdata_72(\time_in|readdata[7]~combout ),
	.readdata_73(\time_out|readdata[7]~q ),
	.readdata_74(\data_o|readdata[7]~q ),
	.readdata_8(\data_i|readdata[8]~combout ),
	.readdata_81(\flags|readdata[8]~q ),
	.readdata_82(\data_o|readdata[8]~q ),
	.readdata_9(\flags|readdata[9]~q ),
	.readdata_10(\flags|readdata[10]~q ),
	.int_nxt_addr_reg_dly_310(\mm_interconnect_0|currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_210(\mm_interconnect_0|currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.int_nxt_addr_reg_dly_311(\mm_interconnect_0|data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_211(\mm_interconnect_0|data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.int_nxt_addr_reg_dly_312(\mm_interconnect_0|tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_212(\mm_interconnect_0|tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.int_nxt_addr_reg_dly_313(\mm_interconnect_0|flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_213(\mm_interconnect_0|flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.int_nxt_addr_reg_dly_314(\mm_interconnect_0|time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_214(\mm_interconnect_0|time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.int_nxt_addr_reg_dly_315(\mm_interconnect_0|tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_215(\mm_interconnect_0|tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.int_nxt_addr_reg_dly_316(\mm_interconnect_0|rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_216(\mm_interconnect_0|rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.clk_clk(\clk_clk~input_o ));

spw_babasu_spw_babasu_pll_0 pll_0(
	.outclk_wire_0(\pll_0|altera_pll_i|outclk_wire[0] ),
	.locked(\pll_0|altera_pll_i|locked_wire[0] ),
	.clk_clk(\clk_clk~input_o ),
	.reset_reset_n(\reset_reset_n~input_o ));

assign \clk_clk~input_o  = clk_clk;

assign \reset_reset_n~input_o  = reset_reset_n;

assign \currentstate_external_connection_export[0]~input_o  = currentstate_external_connection_export[0];

assign \data_o_external_connection_export[0]~input_o  = data_o_external_connection_export[0];

assign \tx_full_external_connection_export~input_o  = tx_full_external_connection_export;

assign \flags_external_connection_export[0]~input_o  = flags_external_connection_export[0];

assign \time_out_external_connection_export[0]~input_o  = time_out_external_connection_export[0];

assign \tick_out_external_connection_export~input_o  = tick_out_external_connection_export;

assign \rx_empty_external_connection_export~input_o  = rx_empty_external_connection_export;

assign \currentstate_external_connection_export[1]~input_o  = currentstate_external_connection_export[1];

assign \time_out_external_connection_export[1]~input_o  = time_out_external_connection_export[1];

assign \data_o_external_connection_export[1]~input_o  = data_o_external_connection_export[1];

assign \flags_external_connection_export[1]~input_o  = flags_external_connection_export[1];

assign \currentstate_external_connection_export[2]~input_o  = currentstate_external_connection_export[2];

assign \time_out_external_connection_export[2]~input_o  = time_out_external_connection_export[2];

assign \data_o_external_connection_export[2]~input_o  = data_o_external_connection_export[2];

assign \flags_external_connection_export[2]~input_o  = flags_external_connection_export[2];

assign \flags_external_connection_export[3]~input_o  = flags_external_connection_export[3];

assign \time_out_external_connection_export[3]~input_o  = time_out_external_connection_export[3];

assign \data_o_external_connection_export[3]~input_o  = data_o_external_connection_export[3];

assign \flags_external_connection_export[4]~input_o  = flags_external_connection_export[4];

assign \time_out_external_connection_export[4]~input_o  = time_out_external_connection_export[4];

assign \data_o_external_connection_export[4]~input_o  = data_o_external_connection_export[4];

assign \flags_external_connection_export[5]~input_o  = flags_external_connection_export[5];

assign \time_out_external_connection_export[5]~input_o  = time_out_external_connection_export[5];

assign \data_o_external_connection_export[5]~input_o  = data_o_external_connection_export[5];

assign \flags_external_connection_export[6]~input_o  = flags_external_connection_export[6];

assign \time_out_external_connection_export[6]~input_o  = time_out_external_connection_export[6];

assign \data_o_external_connection_export[6]~input_o  = data_o_external_connection_export[6];

assign \flags_external_connection_export[7]~input_o  = flags_external_connection_export[7];

assign \time_out_external_connection_export[7]~input_o  = time_out_external_connection_export[7];

assign \data_o_external_connection_export[7]~input_o  = data_o_external_connection_export[7];

assign \flags_external_connection_export[8]~input_o  = flags_external_connection_export[8];

assign \data_o_external_connection_export[8]~input_o  = data_o_external_connection_export[8];

assign \flags_external_connection_export[9]~input_o  = flags_external_connection_export[9];

assign \flags_external_connection_export[10]~input_o  = flags_external_connection_export[10];

assign autostart_external_connection_export = \autostart|data_out~q ;

assign data_i_external_connection_export[0] = \data_i|data_out[0]~q ;

assign data_i_external_connection_export[1] = \data_i|data_out[1]~q ;

assign data_i_external_connection_export[2] = \data_i|data_out[2]~q ;

assign data_i_external_connection_export[3] = \data_i|data_out[3]~q ;

assign data_i_external_connection_export[4] = \data_i|data_out[4]~q ;

assign data_i_external_connection_export[5] = \data_i|data_out[5]~q ;

assign data_i_external_connection_export[6] = \data_i|data_out[6]~q ;

assign data_i_external_connection_export[7] = \data_i|data_out[7]~q ;

assign data_i_external_connection_export[8] = \data_i|data_out[8]~q ;

assign link_disable_external_connection_export = \link_disable|data_out~q ;

assign link_start_external_connection_export = \link_start|data_out~q ;

assign pll_0_locked_export = \pll_0|altera_pll_i|locked_wire[0] ;

assign pll_0_outclk0_clk = \pll_0|altera_pll_i|outclk_wire[0] ;

assign rd_data_external_connection_export = \rd_data|data_out~q ;

assign spill_enable_external_connection_export = \spill_enable|data_out~q ;

assign tick_in_external_connection_export = \tick_in|data_out~q ;

assign time_in_external_connection_export[0] = \time_in|data_out[0]~q ;

assign time_in_external_connection_export[1] = \time_in|data_out[1]~q ;

assign time_in_external_connection_export[2] = \time_in|data_out[2]~q ;

assign time_in_external_connection_export[3] = \time_in|data_out[3]~q ;

assign time_in_external_connection_export[4] = \time_in|data_out[4]~q ;

assign time_in_external_connection_export[5] = \time_in|data_out[5]~q ;

assign time_in_external_connection_export[6] = \time_in|data_out[6]~q ;

assign time_in_external_connection_export[7] = \time_in|data_out[7]~q ;

assign tx_clk_div_external_connection_export[0] = ~ \tx_clk_div|data_out[0]~q ;

assign tx_clk_div_external_connection_export[1] = ~ \tx_clk_div|data_out[1]~q ;

assign tx_clk_div_external_connection_export[2] = \tx_clk_div|data_out[2]~q ;

assign tx_clk_div_external_connection_export[3] = \tx_clk_div|data_out[3]~q ;

assign tx_clk_div_external_connection_export[4] = \tx_clk_div|data_out[4]~q ;

assign tx_clk_div_external_connection_export[5] = \tx_clk_div|data_out[5]~q ;

assign tx_clk_div_external_connection_export[6] = \tx_clk_div|data_out[6]~q ;

assign wr_data_external_connection_export = \wr_data|data_out~q ;

endmodule

module spw_babasu_altera_reset_controller (
	altera_reset_synchronizer_int_chain_out,
	clk_clk,
	reset_reset_n)/* synthesis synthesis_greybox=0 */;
output 	altera_reset_synchronizer_int_chain_out;
input 	clk_clk;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



spw_babasu_altera_reset_synchronizer_3 alt_rst_sync_uq1(
	.altera_reset_synchronizer_int_chain_out1(altera_reset_synchronizer_int_chain_out),
	.clk(clk_clk),
	.reset_reset_n(reset_reset_n));

endmodule

module spw_babasu_altera_reset_controller_1 (
	h2f_rst_n_0,
	altera_reset_synchronizer_int_chain_out,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_rst_n_0;
output 	altera_reset_synchronizer_int_chain_out;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



spw_babasu_altera_reset_synchronizer_1 alt_rst_sync_uq1(
	.h2f_rst_n_0(h2f_rst_n_0),
	.altera_reset_synchronizer_int_chain_out1(altera_reset_synchronizer_int_chain_out),
	.clk(clk_clk));

endmodule

module spw_babasu_altera_reset_synchronizer_1 (
	h2f_rst_n_0,
	altera_reset_synchronizer_int_chain_out1,
	clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_rst_n_0;
output 	altera_reset_synchronizer_int_chain_out1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(h2f_rst_n_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(h2f_rst_n_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(h2f_rst_n_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module spw_babasu_altera_reset_synchronizer_3 (
	altera_reset_synchronizer_int_chain_out1,
	clk,
	reset_reset_n)/* synthesis synthesis_greybox=0 */;
output 	altera_reset_synchronizer_int_chain_out1;
input 	clk;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module spw_babasu_spw_babasu_AUTOSTART (
	data_out1,
	wait_latency_counter_1,
	wait_latency_counter_0,
	m0_write,
	in_data_reg_0,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	reset_n,
	readdata_0,
	clk)/* synthesis synthesis_greybox=0 */;
output 	data_out1;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	m0_write;
input 	in_data_reg_0;
input 	int_nxt_addr_reg_dly_3;
input 	int_nxt_addr_reg_dly_2;
input 	reset_n;
output 	readdata_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always0~0_combout ;
wire \data_out~0_combout ;


dffeas data_out(
	.clk(clk),
	.d(\data_out~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out1),
	.prn(vcc));
defparam data_out.is_wysiwyg = "true";
defparam data_out.power_up = "low";

cyclonev_lcell_comb \readdata[0]~0 (
	.dataa(!data_out1),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[0]~0 .extended_lut = "off";
defparam \readdata[0]~0 .lut_mask = 64'h4040404040404040;
defparam \readdata[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!int_nxt_addr_reg_dly_3),
	.datad(!int_nxt_addr_reg_dly_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'h8000800080008000;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \data_out~0 (
	.dataa(!data_out1),
	.datab(!m0_write),
	.datac(!in_data_reg_0),
	.datad(!\always0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~0 .extended_lut = "off";
defparam \data_out~0 .lut_mask = 64'h5547554755475547;
defparam \data_out~0 .shared_arith = "off";

endmodule

module spw_babasu_spw_babasu_AUTOSTART_1 (
	data_out1,
	wait_latency_counter_1,
	wait_latency_counter_0,
	reset_n,
	m0_write,
	in_data_reg_0,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	readdata_0,
	clk)/* synthesis synthesis_greybox=0 */;
output 	data_out1;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	reset_n;
input 	m0_write;
input 	in_data_reg_0;
input 	int_nxt_addr_reg_dly_3;
input 	int_nxt_addr_reg_dly_2;
output 	readdata_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always0~0_combout ;
wire \data_out~0_combout ;


dffeas data_out(
	.clk(clk),
	.d(\data_out~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out1),
	.prn(vcc));
defparam data_out.is_wysiwyg = "true";
defparam data_out.power_up = "low";

cyclonev_lcell_comb \readdata[0]~0 (
	.dataa(!data_out1),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[0]~0 .extended_lut = "off";
defparam \readdata[0]~0 .lut_mask = 64'h4040404040404040;
defparam \readdata[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!int_nxt_addr_reg_dly_3),
	.datad(!int_nxt_addr_reg_dly_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'h8000800080008000;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \data_out~0 (
	.dataa(!data_out1),
	.datab(!m0_write),
	.datac(!in_data_reg_0),
	.datad(!\always0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~0 .extended_lut = "off";
defparam \data_out~0 .lut_mask = 64'h5547554755475547;
defparam \data_out~0 .shared_arith = "off";

endmodule

module spw_babasu_spw_babasu_AUTOSTART_2 (
	data_out1,
	wait_latency_counter_1,
	wait_latency_counter_0,
	reset_n,
	m0_write,
	in_data_reg_0,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	readdata_0,
	clk)/* synthesis synthesis_greybox=0 */;
output 	data_out1;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	reset_n;
input 	m0_write;
input 	in_data_reg_0;
input 	int_nxt_addr_reg_dly_3;
input 	int_nxt_addr_reg_dly_2;
output 	readdata_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always0~0_combout ;
wire \data_out~0_combout ;


dffeas data_out(
	.clk(clk),
	.d(\data_out~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out1),
	.prn(vcc));
defparam data_out.is_wysiwyg = "true";
defparam data_out.power_up = "low";

cyclonev_lcell_comb \readdata[0]~0 (
	.dataa(!data_out1),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[0]~0 .extended_lut = "off";
defparam \readdata[0]~0 .lut_mask = 64'h4040404040404040;
defparam \readdata[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!int_nxt_addr_reg_dly_3),
	.datad(!int_nxt_addr_reg_dly_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'h8000800080008000;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \data_out~0 (
	.dataa(!data_out1),
	.datab(!m0_write),
	.datac(!in_data_reg_0),
	.datad(!\always0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~0 .extended_lut = "off";
defparam \data_out~0 .lut_mask = 64'h5547554755475547;
defparam \data_out~0 .shared_arith = "off";

endmodule

module spw_babasu_spw_babasu_AUTOSTART_3 (
	data_out1,
	wait_latency_counter_1,
	wait_latency_counter_0,
	reset_n,
	m0_write,
	in_data_reg_0,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	readdata_0,
	clk)/* synthesis synthesis_greybox=0 */;
output 	data_out1;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	reset_n;
input 	m0_write;
input 	in_data_reg_0;
input 	int_nxt_addr_reg_dly_3;
input 	int_nxt_addr_reg_dly_2;
output 	readdata_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always0~0_combout ;
wire \data_out~0_combout ;


dffeas data_out(
	.clk(clk),
	.d(\data_out~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out1),
	.prn(vcc));
defparam data_out.is_wysiwyg = "true";
defparam data_out.power_up = "low";

cyclonev_lcell_comb \readdata[0]~0 (
	.dataa(!data_out1),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[0]~0 .extended_lut = "off";
defparam \readdata[0]~0 .lut_mask = 64'h4040404040404040;
defparam \readdata[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!int_nxt_addr_reg_dly_3),
	.datad(!int_nxt_addr_reg_dly_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'h8000800080008000;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \data_out~0 (
	.dataa(!data_out1),
	.datab(!m0_write),
	.datac(!in_data_reg_0),
	.datad(!\always0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~0 .extended_lut = "off";
defparam \data_out~0 .lut_mask = 64'h5547554755475547;
defparam \data_out~0 .shared_arith = "off";

endmodule

module spw_babasu_spw_babasu_AUTOSTART_4 (
	data_out1,
	wait_latency_counter_1,
	wait_latency_counter_0,
	reset_n,
	m0_write,
	in_data_reg_0,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	readdata_0,
	clk)/* synthesis synthesis_greybox=0 */;
output 	data_out1;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	reset_n;
input 	m0_write;
input 	in_data_reg_0;
input 	int_nxt_addr_reg_dly_3;
input 	int_nxt_addr_reg_dly_2;
output 	readdata_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always0~0_combout ;
wire \data_out~0_combout ;


dffeas data_out(
	.clk(clk),
	.d(\data_out~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out1),
	.prn(vcc));
defparam data_out.is_wysiwyg = "true";
defparam data_out.power_up = "low";

cyclonev_lcell_comb \readdata[0]~0 (
	.dataa(!data_out1),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[0]~0 .extended_lut = "off";
defparam \readdata[0]~0 .lut_mask = 64'h4040404040404040;
defparam \readdata[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!int_nxt_addr_reg_dly_3),
	.datad(!int_nxt_addr_reg_dly_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'h8000800080008000;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \data_out~0 (
	.dataa(!data_out1),
	.datab(!m0_write),
	.datac(!in_data_reg_0),
	.datad(!\always0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~0 .extended_lut = "off";
defparam \data_out~0 .lut_mask = 64'h5547554755475547;
defparam \data_out~0 .shared_arith = "off";

endmodule

module spw_babasu_spw_babasu_AUTOSTART_5 (
	data_out1,
	wait_latency_counter_1,
	wait_latency_counter_0,
	reset_n,
	m0_write,
	in_data_reg_0,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	readdata_0,
	clk)/* synthesis synthesis_greybox=0 */;
output 	data_out1;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	reset_n;
input 	m0_write;
input 	in_data_reg_0;
input 	int_nxt_addr_reg_dly_3;
input 	int_nxt_addr_reg_dly_2;
output 	readdata_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always0~0_combout ;
wire \data_out~0_combout ;


dffeas data_out(
	.clk(clk),
	.d(\data_out~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out1),
	.prn(vcc));
defparam data_out.is_wysiwyg = "true";
defparam data_out.power_up = "low";

cyclonev_lcell_comb \readdata[0]~0 (
	.dataa(!data_out1),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[0]~0 .extended_lut = "off";
defparam \readdata[0]~0 .lut_mask = 64'h4040404040404040;
defparam \readdata[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!int_nxt_addr_reg_dly_3),
	.datad(!int_nxt_addr_reg_dly_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'h8000800080008000;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \data_out~0 (
	.dataa(!data_out1),
	.datab(!m0_write),
	.datac(!in_data_reg_0),
	.datad(!\always0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~0 .extended_lut = "off";
defparam \data_out~0 .lut_mask = 64'h5547554755475547;
defparam \data_out~0 .shared_arith = "off";

endmodule

module spw_babasu_spw_babasu_AUTOSTART_6 (
	data_out1,
	wait_latency_counter_1,
	wait_latency_counter_0,
	reset_n,
	m0_write,
	in_data_reg_0,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	readdata_0,
	clk)/* synthesis synthesis_greybox=0 */;
output 	data_out1;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	reset_n;
input 	m0_write;
input 	in_data_reg_0;
input 	int_nxt_addr_reg_dly_3;
input 	int_nxt_addr_reg_dly_2;
output 	readdata_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always0~0_combout ;
wire \data_out~0_combout ;


dffeas data_out(
	.clk(clk),
	.d(\data_out~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out1),
	.prn(vcc));
defparam data_out.is_wysiwyg = "true";
defparam data_out.power_up = "low";

cyclonev_lcell_comb \readdata[0]~0 (
	.dataa(!data_out1),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[0]~0 .extended_lut = "off";
defparam \readdata[0]~0 .lut_mask = 64'h4040404040404040;
defparam \readdata[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!int_nxt_addr_reg_dly_3),
	.datad(!int_nxt_addr_reg_dly_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'h8000800080008000;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \data_out~0 (
	.dataa(!data_out1),
	.datab(!m0_write),
	.datac(!in_data_reg_0),
	.datad(!\always0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~0 .extended_lut = "off";
defparam \data_out~0 .lut_mask = 64'h5547554755475547;
defparam \data_out~0 .shared_arith = "off";

endmodule

module spw_babasu_spw_babasu_CURRENTSTATE (
	altera_reset_synchronizer_int_chain_out,
	readdata_0,
	readdata_1,
	readdata_2,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	clk_clk,
	currentstate_external_connection_export_0,
	currentstate_external_connection_export_1,
	currentstate_external_connection_export_2)/* synthesis synthesis_greybox=0 */;
input 	altera_reset_synchronizer_int_chain_out;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
input 	int_nxt_addr_reg_dly_3;
input 	int_nxt_addr_reg_dly_2;
input 	clk_clk;
input 	currentstate_external_connection_export_0;
input 	currentstate_external_connection_export_1;
input 	currentstate_external_connection_export_2;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_mux_out[0]~0_combout ;
wire \read_mux_out[1]~1_combout ;
wire \read_mux_out[2]~2_combout ;


dffeas \readdata[0] (
	.clk(clk_clk),
	.d(\read_mux_out[0]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

dffeas \readdata[1] (
	.clk(clk_clk),
	.d(\read_mux_out[1]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_1),
	.prn(vcc));
defparam \readdata[1] .is_wysiwyg = "true";
defparam \readdata[1] .power_up = "low";

dffeas \readdata[2] (
	.clk(clk_clk),
	.d(\read_mux_out[2]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_2),
	.prn(vcc));
defparam \readdata[2] .is_wysiwyg = "true";
defparam \readdata[2] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[0]~0 (
	.dataa(!currentstate_external_connection_export_0),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[0]~0 .extended_lut = "off";
defparam \read_mux_out[0]~0 .lut_mask = 64'h4040404040404040;
defparam \read_mux_out[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[1]~1 (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!currentstate_external_connection_export_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[1]~1 .extended_lut = "off";
defparam \read_mux_out[1]~1 .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[2]~2 (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!currentstate_external_connection_export_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[2]~2 .extended_lut = "off";
defparam \read_mux_out[2]~2 .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[2]~2 .shared_arith = "off";

endmodule

module spw_babasu_spw_babasu_DATA_I (
	data_out_0,
	data_out_1,
	data_out_2,
	data_out_3,
	data_out_4,
	data_out_5,
	data_out_6,
	data_out_7,
	data_out_8,
	wait_latency_counter_1,
	wait_latency_counter_0,
	reset_n,
	writedata,
	m0_write,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	readdata_4,
	readdata_5,
	readdata_6,
	readdata_7,
	readdata_8,
	clk)/* synthesis synthesis_greybox=0 */;
output 	data_out_0;
output 	data_out_1;
output 	data_out_2;
output 	data_out_3;
output 	data_out_4;
output 	data_out_5;
output 	data_out_6;
output 	data_out_7;
output 	data_out_8;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	reset_n;
input 	[31:0] writedata;
input 	m0_write;
input 	int_nxt_addr_reg_dly_3;
input 	int_nxt_addr_reg_dly_2;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
output 	readdata_4;
output 	readdata_5;
output 	readdata_6;
output 	readdata_7;
output 	readdata_8;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always0~0_combout ;


dffeas \data_out[0] (
	.clk(clk),
	.d(writedata[0]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_0),
	.prn(vcc));
defparam \data_out[0] .is_wysiwyg = "true";
defparam \data_out[0] .power_up = "low";

dffeas \data_out[1] (
	.clk(clk),
	.d(writedata[1]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_1),
	.prn(vcc));
defparam \data_out[1] .is_wysiwyg = "true";
defparam \data_out[1] .power_up = "low";

dffeas \data_out[2] (
	.clk(clk),
	.d(writedata[2]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_2),
	.prn(vcc));
defparam \data_out[2] .is_wysiwyg = "true";
defparam \data_out[2] .power_up = "low";

dffeas \data_out[3] (
	.clk(clk),
	.d(writedata[3]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_3),
	.prn(vcc));
defparam \data_out[3] .is_wysiwyg = "true";
defparam \data_out[3] .power_up = "low";

dffeas \data_out[4] (
	.clk(clk),
	.d(writedata[4]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_4),
	.prn(vcc));
defparam \data_out[4] .is_wysiwyg = "true";
defparam \data_out[4] .power_up = "low";

dffeas \data_out[5] (
	.clk(clk),
	.d(writedata[5]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_5),
	.prn(vcc));
defparam \data_out[5] .is_wysiwyg = "true";
defparam \data_out[5] .power_up = "low";

dffeas \data_out[6] (
	.clk(clk),
	.d(writedata[6]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_6),
	.prn(vcc));
defparam \data_out[6] .is_wysiwyg = "true";
defparam \data_out[6] .power_up = "low";

dffeas \data_out[7] (
	.clk(clk),
	.d(writedata[7]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_7),
	.prn(vcc));
defparam \data_out[7] .is_wysiwyg = "true";
defparam \data_out[7] .power_up = "low";

dffeas \data_out[8] (
	.clk(clk),
	.d(writedata[8]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_8),
	.prn(vcc));
defparam \data_out[8] .is_wysiwyg = "true";
defparam \data_out[8] .power_up = "low";

cyclonev_lcell_comb \readdata[0] (
	.dataa(!data_out_0),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[0] .extended_lut = "off";
defparam \readdata[0] .lut_mask = 64'h4040404040404040;
defparam \readdata[0] .shared_arith = "off";

cyclonev_lcell_comb \readdata[1] (
	.dataa(!data_out_1),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[1] .extended_lut = "off";
defparam \readdata[1] .lut_mask = 64'h4040404040404040;
defparam \readdata[1] .shared_arith = "off";

cyclonev_lcell_comb \readdata[2] (
	.dataa(!data_out_2),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[2] .extended_lut = "off";
defparam \readdata[2] .lut_mask = 64'h4040404040404040;
defparam \readdata[2] .shared_arith = "off";

cyclonev_lcell_comb \readdata[3] (
	.dataa(!data_out_3),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[3] .extended_lut = "off";
defparam \readdata[3] .lut_mask = 64'h4040404040404040;
defparam \readdata[3] .shared_arith = "off";

cyclonev_lcell_comb \readdata[4] (
	.dataa(!data_out_4),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[4] .extended_lut = "off";
defparam \readdata[4] .lut_mask = 64'h4040404040404040;
defparam \readdata[4] .shared_arith = "off";

cyclonev_lcell_comb \readdata[5] (
	.dataa(!data_out_5),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[5] .extended_lut = "off";
defparam \readdata[5] .lut_mask = 64'h4040404040404040;
defparam \readdata[5] .shared_arith = "off";

cyclonev_lcell_comb \readdata[6] (
	.dataa(!data_out_6),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_6),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[6] .extended_lut = "off";
defparam \readdata[6] .lut_mask = 64'h4040404040404040;
defparam \readdata[6] .shared_arith = "off";

cyclonev_lcell_comb \readdata[7] (
	.dataa(!data_out_7),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_7),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[7] .extended_lut = "off";
defparam \readdata[7] .lut_mask = 64'h4040404040404040;
defparam \readdata[7] .shared_arith = "off";

cyclonev_lcell_comb \readdata[8] (
	.dataa(!data_out_8),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[8] .extended_lut = "off";
defparam \readdata[8] .lut_mask = 64'h4040404040404040;
defparam \readdata[8] .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!m0_write),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(!int_nxt_addr_reg_dly_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'h0800000008000000;
defparam \always0~0 .shared_arith = "off";

endmodule

module spw_babasu_spw_babasu_DATA_O (
	altera_reset_synchronizer_int_chain_out,
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	readdata_4,
	readdata_5,
	readdata_6,
	readdata_7,
	readdata_8,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	clk_clk,
	data_o_external_connection_export_0,
	data_o_external_connection_export_1,
	data_o_external_connection_export_2,
	data_o_external_connection_export_3,
	data_o_external_connection_export_4,
	data_o_external_connection_export_5,
	data_o_external_connection_export_6,
	data_o_external_connection_export_7,
	data_o_external_connection_export_8)/* synthesis synthesis_greybox=0 */;
input 	altera_reset_synchronizer_int_chain_out;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
output 	readdata_4;
output 	readdata_5;
output 	readdata_6;
output 	readdata_7;
output 	readdata_8;
input 	int_nxt_addr_reg_dly_3;
input 	int_nxt_addr_reg_dly_2;
input 	clk_clk;
input 	data_o_external_connection_export_0;
input 	data_o_external_connection_export_1;
input 	data_o_external_connection_export_2;
input 	data_o_external_connection_export_3;
input 	data_o_external_connection_export_4;
input 	data_o_external_connection_export_5;
input 	data_o_external_connection_export_6;
input 	data_o_external_connection_export_7;
input 	data_o_external_connection_export_8;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_mux_out[0]~combout ;
wire \read_mux_out[1]~combout ;
wire \read_mux_out[2]~combout ;
wire \read_mux_out[3]~combout ;
wire \read_mux_out[4]~combout ;
wire \read_mux_out[5]~combout ;
wire \read_mux_out[6]~combout ;
wire \read_mux_out[7]~combout ;
wire \read_mux_out[8]~combout ;


dffeas \readdata[0] (
	.clk(clk_clk),
	.d(\read_mux_out[0]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

dffeas \readdata[1] (
	.clk(clk_clk),
	.d(\read_mux_out[1]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_1),
	.prn(vcc));
defparam \readdata[1] .is_wysiwyg = "true";
defparam \readdata[1] .power_up = "low";

dffeas \readdata[2] (
	.clk(clk_clk),
	.d(\read_mux_out[2]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_2),
	.prn(vcc));
defparam \readdata[2] .is_wysiwyg = "true";
defparam \readdata[2] .power_up = "low";

dffeas \readdata[3] (
	.clk(clk_clk),
	.d(\read_mux_out[3]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_3),
	.prn(vcc));
defparam \readdata[3] .is_wysiwyg = "true";
defparam \readdata[3] .power_up = "low";

dffeas \readdata[4] (
	.clk(clk_clk),
	.d(\read_mux_out[4]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_4),
	.prn(vcc));
defparam \readdata[4] .is_wysiwyg = "true";
defparam \readdata[4] .power_up = "low";

dffeas \readdata[5] (
	.clk(clk_clk),
	.d(\read_mux_out[5]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_5),
	.prn(vcc));
defparam \readdata[5] .is_wysiwyg = "true";
defparam \readdata[5] .power_up = "low";

dffeas \readdata[6] (
	.clk(clk_clk),
	.d(\read_mux_out[6]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_6),
	.prn(vcc));
defparam \readdata[6] .is_wysiwyg = "true";
defparam \readdata[6] .power_up = "low";

dffeas \readdata[7] (
	.clk(clk_clk),
	.d(\read_mux_out[7]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_7),
	.prn(vcc));
defparam \readdata[7] .is_wysiwyg = "true";
defparam \readdata[7] .power_up = "low";

dffeas \readdata[8] (
	.clk(clk_clk),
	.d(\read_mux_out[8]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_8),
	.prn(vcc));
defparam \readdata[8] .is_wysiwyg = "true";
defparam \readdata[8] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[0] (
	.dataa(!data_o_external_connection_export_0),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[0] .extended_lut = "off";
defparam \read_mux_out[0] .lut_mask = 64'h4040404040404040;
defparam \read_mux_out[0] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[1] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!data_o_external_connection_export_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[1] .extended_lut = "off";
defparam \read_mux_out[1] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[1] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[2] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!data_o_external_connection_export_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[2] .extended_lut = "off";
defparam \read_mux_out[2] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[2] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[3] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!data_o_external_connection_export_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[3] .extended_lut = "off";
defparam \read_mux_out[3] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[3] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[4] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!data_o_external_connection_export_4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[4]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[4] .extended_lut = "off";
defparam \read_mux_out[4] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[4] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[5] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!data_o_external_connection_export_5),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[5]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[5] .extended_lut = "off";
defparam \read_mux_out[5] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[5] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[6] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!data_o_external_connection_export_6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[6]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[6] .extended_lut = "off";
defparam \read_mux_out[6] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[6] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[7] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!data_o_external_connection_export_7),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[7]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[7] .extended_lut = "off";
defparam \read_mux_out[7] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[7] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[8] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!data_o_external_connection_export_8),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[8]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[8] .extended_lut = "off";
defparam \read_mux_out[8] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[8] .shared_arith = "off";

endmodule

module spw_babasu_spw_babasu_FLAGS (
	altera_reset_synchronizer_int_chain_out,
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	readdata_4,
	readdata_5,
	readdata_6,
	readdata_7,
	readdata_8,
	readdata_9,
	readdata_10,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	clk_clk,
	flags_external_connection_export_0,
	flags_external_connection_export_1,
	flags_external_connection_export_2,
	flags_external_connection_export_3,
	flags_external_connection_export_4,
	flags_external_connection_export_5,
	flags_external_connection_export_6,
	flags_external_connection_export_7,
	flags_external_connection_export_8,
	flags_external_connection_export_9,
	flags_external_connection_export_10)/* synthesis synthesis_greybox=0 */;
input 	altera_reset_synchronizer_int_chain_out;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
output 	readdata_4;
output 	readdata_5;
output 	readdata_6;
output 	readdata_7;
output 	readdata_8;
output 	readdata_9;
output 	readdata_10;
input 	int_nxt_addr_reg_dly_3;
input 	int_nxt_addr_reg_dly_2;
input 	clk_clk;
input 	flags_external_connection_export_0;
input 	flags_external_connection_export_1;
input 	flags_external_connection_export_2;
input 	flags_external_connection_export_3;
input 	flags_external_connection_export_4;
input 	flags_external_connection_export_5;
input 	flags_external_connection_export_6;
input 	flags_external_connection_export_7;
input 	flags_external_connection_export_8;
input 	flags_external_connection_export_9;
input 	flags_external_connection_export_10;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_mux_out[0]~combout ;
wire \read_mux_out[1]~combout ;
wire \read_mux_out[2]~combout ;
wire \read_mux_out[3]~combout ;
wire \read_mux_out[4]~combout ;
wire \read_mux_out[5]~combout ;
wire \read_mux_out[6]~combout ;
wire \read_mux_out[7]~combout ;
wire \read_mux_out[8]~combout ;
wire \read_mux_out[9]~combout ;
wire \read_mux_out[10]~combout ;


dffeas \readdata[0] (
	.clk(clk_clk),
	.d(\read_mux_out[0]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

dffeas \readdata[1] (
	.clk(clk_clk),
	.d(\read_mux_out[1]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_1),
	.prn(vcc));
defparam \readdata[1] .is_wysiwyg = "true";
defparam \readdata[1] .power_up = "low";

dffeas \readdata[2] (
	.clk(clk_clk),
	.d(\read_mux_out[2]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_2),
	.prn(vcc));
defparam \readdata[2] .is_wysiwyg = "true";
defparam \readdata[2] .power_up = "low";

dffeas \readdata[3] (
	.clk(clk_clk),
	.d(\read_mux_out[3]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_3),
	.prn(vcc));
defparam \readdata[3] .is_wysiwyg = "true";
defparam \readdata[3] .power_up = "low";

dffeas \readdata[4] (
	.clk(clk_clk),
	.d(\read_mux_out[4]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_4),
	.prn(vcc));
defparam \readdata[4] .is_wysiwyg = "true";
defparam \readdata[4] .power_up = "low";

dffeas \readdata[5] (
	.clk(clk_clk),
	.d(\read_mux_out[5]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_5),
	.prn(vcc));
defparam \readdata[5] .is_wysiwyg = "true";
defparam \readdata[5] .power_up = "low";

dffeas \readdata[6] (
	.clk(clk_clk),
	.d(\read_mux_out[6]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_6),
	.prn(vcc));
defparam \readdata[6] .is_wysiwyg = "true";
defparam \readdata[6] .power_up = "low";

dffeas \readdata[7] (
	.clk(clk_clk),
	.d(\read_mux_out[7]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_7),
	.prn(vcc));
defparam \readdata[7] .is_wysiwyg = "true";
defparam \readdata[7] .power_up = "low";

dffeas \readdata[8] (
	.clk(clk_clk),
	.d(\read_mux_out[8]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_8),
	.prn(vcc));
defparam \readdata[8] .is_wysiwyg = "true";
defparam \readdata[8] .power_up = "low";

dffeas \readdata[9] (
	.clk(clk_clk),
	.d(\read_mux_out[9]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_9),
	.prn(vcc));
defparam \readdata[9] .is_wysiwyg = "true";
defparam \readdata[9] .power_up = "low";

dffeas \readdata[10] (
	.clk(clk_clk),
	.d(\read_mux_out[10]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_10),
	.prn(vcc));
defparam \readdata[10] .is_wysiwyg = "true";
defparam \readdata[10] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[0] (
	.dataa(!flags_external_connection_export_0),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[0] .extended_lut = "off";
defparam \read_mux_out[0] .lut_mask = 64'h4040404040404040;
defparam \read_mux_out[0] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[1] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!flags_external_connection_export_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[1] .extended_lut = "off";
defparam \read_mux_out[1] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[1] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[2] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!flags_external_connection_export_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[2] .extended_lut = "off";
defparam \read_mux_out[2] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[2] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[3] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!flags_external_connection_export_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[3] .extended_lut = "off";
defparam \read_mux_out[3] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[3] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[4] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!flags_external_connection_export_4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[4]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[4] .extended_lut = "off";
defparam \read_mux_out[4] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[4] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[5] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!flags_external_connection_export_5),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[5]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[5] .extended_lut = "off";
defparam \read_mux_out[5] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[5] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[6] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!flags_external_connection_export_6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[6]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[6] .extended_lut = "off";
defparam \read_mux_out[6] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[6] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[7] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!flags_external_connection_export_7),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[7]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[7] .extended_lut = "off";
defparam \read_mux_out[7] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[7] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[8] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!flags_external_connection_export_8),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[8]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[8] .extended_lut = "off";
defparam \read_mux_out[8] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[8] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[9] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!flags_external_connection_export_9),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[9]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[9] .extended_lut = "off";
defparam \read_mux_out[9] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[9] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[10] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!flags_external_connection_export_10),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[10]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[10] .extended_lut = "off";
defparam \read_mux_out[10] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[10] .shared_arith = "off";

endmodule

module spw_babasu_spw_babasu_hps_0 (
	h2f_rst_n_0,
	h2f_ARVALID_0,
	h2f_AWVALID_0,
	h2f_BREADY_0,
	h2f_RREADY_0,
	h2f_WLAST_0,
	h2f_WVALID_0,
	h2f_ARADDR_0,
	h2f_ARADDR_1,
	h2f_ARADDR_2,
	h2f_ARADDR_3,
	h2f_ARADDR_4,
	h2f_ARADDR_5,
	h2f_ARADDR_6,
	h2f_ARADDR_7,
	h2f_ARADDR_8,
	h2f_ARBURST_0,
	h2f_ARBURST_1,
	h2f_ARID_0,
	h2f_ARID_1,
	h2f_ARID_2,
	h2f_ARID_3,
	h2f_ARID_4,
	h2f_ARID_5,
	h2f_ARID_6,
	h2f_ARID_7,
	h2f_ARID_8,
	h2f_ARID_9,
	h2f_ARID_10,
	h2f_ARID_11,
	h2f_ARLEN_0,
	h2f_ARLEN_1,
	h2f_ARLEN_2,
	h2f_ARLEN_3,
	h2f_ARSIZE_0,
	h2f_ARSIZE_1,
	h2f_ARSIZE_2,
	h2f_AWADDR_0,
	h2f_AWADDR_1,
	h2f_AWADDR_2,
	h2f_AWADDR_3,
	h2f_AWADDR_4,
	h2f_AWADDR_5,
	h2f_AWADDR_6,
	h2f_AWADDR_7,
	h2f_AWADDR_8,
	h2f_AWBURST_0,
	h2f_AWBURST_1,
	h2f_AWID_0,
	h2f_AWID_1,
	h2f_AWID_2,
	h2f_AWID_3,
	h2f_AWID_4,
	h2f_AWID_5,
	h2f_AWID_6,
	h2f_AWID_7,
	h2f_AWID_8,
	h2f_AWID_9,
	h2f_AWID_10,
	h2f_AWID_11,
	h2f_AWLEN_0,
	h2f_AWLEN_1,
	h2f_AWLEN_2,
	h2f_AWLEN_3,
	h2f_AWSIZE_0,
	h2f_AWSIZE_1,
	h2f_AWSIZE_2,
	h2f_WDATA_0,
	h2f_WDATA_1,
	h2f_WDATA_2,
	h2f_WDATA_3,
	h2f_WDATA_4,
	h2f_WDATA_5,
	h2f_WDATA_6,
	h2f_WDATA_7,
	h2f_WDATA_8,
	h2f_WSTRB_0,
	h2f_WSTRB_1,
	h2f_WSTRB_2,
	h2f_WSTRB_3,
	cmd_sink_ready,
	nonposted_cmd_accepted,
	WideOr1,
	src_payload_0,
	WideOr11,
	nonposted_cmd_accepted1,
	src_data_105,
	src_data_106,
	src_data_107,
	src_data_108,
	src_data_109,
	src_data_110,
	src_data_111,
	src_data_112,
	src_data_113,
	src_data_114,
	src_data_115,
	src_data_116,
	src_data_0,
	src_payload,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_data_1051,
	src_data_1061,
	src_data_1071,
	src_data_1081,
	src_data_1091,
	src_data_1101,
	src_data_1111,
	src_data_1121,
	src_data_1131,
	src_data_1141,
	src_data_1151,
	src_data_1161,
	clk_clk)/* synthesis synthesis_greybox=0 */;
output 	h2f_rst_n_0;
output 	h2f_ARVALID_0;
output 	h2f_AWVALID_0;
output 	h2f_BREADY_0;
output 	h2f_RREADY_0;
output 	h2f_WLAST_0;
output 	h2f_WVALID_0;
output 	h2f_ARADDR_0;
output 	h2f_ARADDR_1;
output 	h2f_ARADDR_2;
output 	h2f_ARADDR_3;
output 	h2f_ARADDR_4;
output 	h2f_ARADDR_5;
output 	h2f_ARADDR_6;
output 	h2f_ARADDR_7;
output 	h2f_ARADDR_8;
output 	h2f_ARBURST_0;
output 	h2f_ARBURST_1;
output 	h2f_ARID_0;
output 	h2f_ARID_1;
output 	h2f_ARID_2;
output 	h2f_ARID_3;
output 	h2f_ARID_4;
output 	h2f_ARID_5;
output 	h2f_ARID_6;
output 	h2f_ARID_7;
output 	h2f_ARID_8;
output 	h2f_ARID_9;
output 	h2f_ARID_10;
output 	h2f_ARID_11;
output 	h2f_ARLEN_0;
output 	h2f_ARLEN_1;
output 	h2f_ARLEN_2;
output 	h2f_ARLEN_3;
output 	h2f_ARSIZE_0;
output 	h2f_ARSIZE_1;
output 	h2f_ARSIZE_2;
output 	h2f_AWADDR_0;
output 	h2f_AWADDR_1;
output 	h2f_AWADDR_2;
output 	h2f_AWADDR_3;
output 	h2f_AWADDR_4;
output 	h2f_AWADDR_5;
output 	h2f_AWADDR_6;
output 	h2f_AWADDR_7;
output 	h2f_AWADDR_8;
output 	h2f_AWBURST_0;
output 	h2f_AWBURST_1;
output 	h2f_AWID_0;
output 	h2f_AWID_1;
output 	h2f_AWID_2;
output 	h2f_AWID_3;
output 	h2f_AWID_4;
output 	h2f_AWID_5;
output 	h2f_AWID_6;
output 	h2f_AWID_7;
output 	h2f_AWID_8;
output 	h2f_AWID_9;
output 	h2f_AWID_10;
output 	h2f_AWID_11;
output 	h2f_AWLEN_0;
output 	h2f_AWLEN_1;
output 	h2f_AWLEN_2;
output 	h2f_AWLEN_3;
output 	h2f_AWSIZE_0;
output 	h2f_AWSIZE_1;
output 	h2f_AWSIZE_2;
output 	h2f_WDATA_0;
output 	h2f_WDATA_1;
output 	h2f_WDATA_2;
output 	h2f_WDATA_3;
output 	h2f_WDATA_4;
output 	h2f_WDATA_5;
output 	h2f_WDATA_6;
output 	h2f_WDATA_7;
output 	h2f_WDATA_8;
output 	h2f_WSTRB_0;
output 	h2f_WSTRB_1;
output 	h2f_WSTRB_2;
output 	h2f_WSTRB_3;
input 	cmd_sink_ready;
input 	nonposted_cmd_accepted;
input 	WideOr1;
input 	src_payload_0;
input 	WideOr11;
input 	nonposted_cmd_accepted1;
input 	src_data_105;
input 	src_data_106;
input 	src_data_107;
input 	src_data_108;
input 	src_data_109;
input 	src_data_110;
input 	src_data_111;
input 	src_data_112;
input 	src_data_113;
input 	src_data_114;
input 	src_data_115;
input 	src_data_116;
input 	src_data_0;
input 	src_payload;
input 	src_payload1;
input 	src_payload2;
input 	src_payload3;
input 	src_payload4;
input 	src_payload5;
input 	src_payload6;
input 	src_payload7;
input 	src_payload8;
input 	src_payload9;
input 	src_data_1051;
input 	src_data_1061;
input 	src_data_1071;
input 	src_data_1081;
input 	src_data_1091;
input 	src_data_1101;
input 	src_data_1111;
input 	src_data_1121;
input 	src_data_1131;
input 	src_data_1141;
input 	src_data_1151;
input 	src_data_1161;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



spw_babasu_spw_babasu_hps_0_fpga_interfaces fpga_interfaces(
	.h2f_rst_n({h2f_rst_n_0}),
	.h2f_ARVALID({h2f_ARVALID_0}),
	.h2f_AWVALID({h2f_AWVALID_0}),
	.h2f_BREADY({h2f_BREADY_0}),
	.h2f_RREADY({h2f_RREADY_0}),
	.h2f_WLAST({h2f_WLAST_0}),
	.h2f_WVALID({h2f_WVALID_0}),
	.h2f_ARADDR({h2f_ARADDR_unconnected_wire_29,h2f_ARADDR_unconnected_wire_28,h2f_ARADDR_unconnected_wire_27,h2f_ARADDR_unconnected_wire_26,h2f_ARADDR_unconnected_wire_25,h2f_ARADDR_unconnected_wire_24,h2f_ARADDR_unconnected_wire_23,h2f_ARADDR_unconnected_wire_22,
h2f_ARADDR_unconnected_wire_21,h2f_ARADDR_unconnected_wire_20,h2f_ARADDR_unconnected_wire_19,h2f_ARADDR_unconnected_wire_18,h2f_ARADDR_unconnected_wire_17,h2f_ARADDR_unconnected_wire_16,h2f_ARADDR_unconnected_wire_15,h2f_ARADDR_unconnected_wire_14,
h2f_ARADDR_unconnected_wire_13,h2f_ARADDR_unconnected_wire_12,h2f_ARADDR_unconnected_wire_11,h2f_ARADDR_unconnected_wire_10,h2f_ARADDR_unconnected_wire_9,h2f_ARADDR_8,h2f_ARADDR_7,h2f_ARADDR_6,h2f_ARADDR_5,h2f_ARADDR_4,h2f_ARADDR_3,h2f_ARADDR_2,h2f_ARADDR_1,
h2f_ARADDR_0}),
	.h2f_ARBURST({h2f_ARBURST_1,h2f_ARBURST_0}),
	.h2f_ARID({h2f_ARID_11,h2f_ARID_10,h2f_ARID_9,h2f_ARID_8,h2f_ARID_7,h2f_ARID_6,h2f_ARID_5,h2f_ARID_4,h2f_ARID_3,h2f_ARID_2,h2f_ARID_1,h2f_ARID_0}),
	.h2f_ARLEN({h2f_ARLEN_3,h2f_ARLEN_2,h2f_ARLEN_1,h2f_ARLEN_0}),
	.h2f_ARSIZE({h2f_ARSIZE_2,h2f_ARSIZE_1,h2f_ARSIZE_0}),
	.h2f_AWADDR({h2f_AWADDR_unconnected_wire_29,h2f_AWADDR_unconnected_wire_28,h2f_AWADDR_unconnected_wire_27,h2f_AWADDR_unconnected_wire_26,h2f_AWADDR_unconnected_wire_25,h2f_AWADDR_unconnected_wire_24,h2f_AWADDR_unconnected_wire_23,h2f_AWADDR_unconnected_wire_22,
h2f_AWADDR_unconnected_wire_21,h2f_AWADDR_unconnected_wire_20,h2f_AWADDR_unconnected_wire_19,h2f_AWADDR_unconnected_wire_18,h2f_AWADDR_unconnected_wire_17,h2f_AWADDR_unconnected_wire_16,h2f_AWADDR_unconnected_wire_15,h2f_AWADDR_unconnected_wire_14,
h2f_AWADDR_unconnected_wire_13,h2f_AWADDR_unconnected_wire_12,h2f_AWADDR_unconnected_wire_11,h2f_AWADDR_unconnected_wire_10,h2f_AWADDR_unconnected_wire_9,h2f_AWADDR_8,h2f_AWADDR_7,h2f_AWADDR_6,h2f_AWADDR_5,h2f_AWADDR_4,h2f_AWADDR_3,h2f_AWADDR_2,h2f_AWADDR_1,
h2f_AWADDR_0}),
	.h2f_AWBURST({h2f_AWBURST_1,h2f_AWBURST_0}),
	.h2f_AWID({h2f_AWID_11,h2f_AWID_10,h2f_AWID_9,h2f_AWID_8,h2f_AWID_7,h2f_AWID_6,h2f_AWID_5,h2f_AWID_4,h2f_AWID_3,h2f_AWID_2,h2f_AWID_1,h2f_AWID_0}),
	.h2f_AWLEN({h2f_AWLEN_3,h2f_AWLEN_2,h2f_AWLEN_1,h2f_AWLEN_0}),
	.h2f_AWSIZE({h2f_AWSIZE_2,h2f_AWSIZE_1,h2f_AWSIZE_0}),
	.h2f_WDATA({h2f_WDATA_unconnected_wire_31,h2f_WDATA_unconnected_wire_30,h2f_WDATA_unconnected_wire_29,h2f_WDATA_unconnected_wire_28,h2f_WDATA_unconnected_wire_27,h2f_WDATA_unconnected_wire_26,h2f_WDATA_unconnected_wire_25,h2f_WDATA_unconnected_wire_24,
h2f_WDATA_unconnected_wire_23,h2f_WDATA_unconnected_wire_22,h2f_WDATA_unconnected_wire_21,h2f_WDATA_unconnected_wire_20,h2f_WDATA_unconnected_wire_19,h2f_WDATA_unconnected_wire_18,h2f_WDATA_unconnected_wire_17,h2f_WDATA_unconnected_wire_16,
h2f_WDATA_unconnected_wire_15,h2f_WDATA_unconnected_wire_14,h2f_WDATA_unconnected_wire_13,h2f_WDATA_unconnected_wire_12,h2f_WDATA_unconnected_wire_11,h2f_WDATA_unconnected_wire_10,h2f_WDATA_unconnected_wire_9,h2f_WDATA_8,h2f_WDATA_7,h2f_WDATA_6,h2f_WDATA_5,
h2f_WDATA_4,h2f_WDATA_3,h2f_WDATA_2,h2f_WDATA_1,h2f_WDATA_0}),
	.h2f_WSTRB({h2f_WSTRB_3,h2f_WSTRB_2,h2f_WSTRB_1,h2f_WSTRB_0}),
	.h2f_ARREADY({cmd_sink_ready}),
	.h2f_AWREADY({nonposted_cmd_accepted}),
	.h2f_BVALID({WideOr1}),
	.h2f_RLAST({src_payload_0}),
	.h2f_RVALID({WideOr11}),
	.h2f_WREADY({nonposted_cmd_accepted1}),
	.h2f_BID({src_data_116,src_data_115,src_data_114,src_data_113,src_data_112,src_data_111,src_data_110,src_data_109,src_data_108,src_data_107,src_data_106,src_data_105}),
	.h2f_RDATA({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_payload9,src_payload8,src_payload7,src_payload6,src_payload5,src_payload4,src_payload3,src_payload2,src_payload1,src_payload,src_data_0}),
	.h2f_RID({src_data_1161,src_data_1151,src_data_1141,src_data_1131,src_data_1121,src_data_1111,src_data_1101,src_data_1091,src_data_1081,src_data_1071,src_data_1061,src_data_1051}),
	.h2f_axi_clk({clk_clk}));

endmodule

module spw_babasu_spw_babasu_hps_0_fpga_interfaces (
	h2f_rst_n,
	h2f_ARVALID,
	h2f_AWVALID,
	h2f_BREADY,
	h2f_RREADY,
	h2f_WLAST,
	h2f_WVALID,
	h2f_ARADDR,
	h2f_ARBURST,
	h2f_ARID,
	h2f_ARLEN,
	h2f_ARSIZE,
	h2f_AWADDR,
	h2f_AWBURST,
	h2f_AWID,
	h2f_AWLEN,
	h2f_AWSIZE,
	h2f_WDATA,
	h2f_WSTRB,
	h2f_ARREADY,
	h2f_AWREADY,
	h2f_BVALID,
	h2f_RLAST,
	h2f_RVALID,
	h2f_WREADY,
	h2f_BID,
	h2f_RDATA,
	h2f_RID,
	h2f_axi_clk)/* synthesis synthesis_greybox=0 */;
output 	[0:0] h2f_rst_n;
output 	[0:0] h2f_ARVALID;
output 	[0:0] h2f_AWVALID;
output 	[0:0] h2f_BREADY;
output 	[0:0] h2f_RREADY;
output 	[0:0] h2f_WLAST;
output 	[0:0] h2f_WVALID;
output 	[29:0] h2f_ARADDR;
output 	[1:0] h2f_ARBURST;
output 	[11:0] h2f_ARID;
output 	[3:0] h2f_ARLEN;
output 	[2:0] h2f_ARSIZE;
output 	[29:0] h2f_AWADDR;
output 	[1:0] h2f_AWBURST;
output 	[11:0] h2f_AWID;
output 	[3:0] h2f_AWLEN;
output 	[2:0] h2f_AWSIZE;
output 	[31:0] h2f_WDATA;
output 	[3:0] h2f_WSTRB;
input 	[0:0] h2f_ARREADY;
input 	[0:0] h2f_AWREADY;
input 	[0:0] h2f_BVALID;
input 	[0:0] h2f_RLAST;
input 	[0:0] h2f_RVALID;
input 	[0:0] h2f_WREADY;
input 	[11:0] h2f_BID;
input 	[31:0] h2f_RDATA;
input 	[11:0] h2f_RID;
input 	[0:0] h2f_axi_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \debug_apb~O_P_ADDR_31 ;
wire \tpiu~trace_data ;
wire \tpiu~O_TRACE_DATA1 ;
wire \tpiu~O_TRACE_DATA2 ;
wire \tpiu~O_TRACE_DATA3 ;
wire \tpiu~O_TRACE_DATA4 ;
wire \tpiu~O_TRACE_DATA5 ;
wire \tpiu~O_TRACE_DATA6 ;
wire \tpiu~O_TRACE_DATA7 ;
wire \tpiu~O_TRACE_DATA8 ;
wire \tpiu~O_TRACE_DATA9 ;
wire \tpiu~O_TRACE_DATA10 ;
wire \tpiu~O_TRACE_DATA11 ;
wire \tpiu~O_TRACE_DATA12 ;
wire \tpiu~O_TRACE_DATA13 ;
wire \tpiu~O_TRACE_DATA14 ;
wire \tpiu~O_TRACE_DATA15 ;
wire \tpiu~O_TRACE_DATA16 ;
wire \tpiu~O_TRACE_DATA17 ;
wire \tpiu~O_TRACE_DATA18 ;
wire \tpiu~O_TRACE_DATA19 ;
wire \tpiu~O_TRACE_DATA20 ;
wire \tpiu~O_TRACE_DATA21 ;
wire \tpiu~O_TRACE_DATA22 ;
wire \tpiu~O_TRACE_DATA23 ;
wire \tpiu~O_TRACE_DATA24 ;
wire \tpiu~O_TRACE_DATA25 ;
wire \tpiu~O_TRACE_DATA26 ;
wire \tpiu~O_TRACE_DATA27 ;
wire \tpiu~O_TRACE_DATA28 ;
wire \tpiu~O_TRACE_DATA29 ;
wire \tpiu~O_TRACE_DATA30 ;
wire \tpiu~O_TRACE_DATA31 ;
wire \boot_from_fpga~fake_dout ;
wire \fpga2hps~arready ;
wire \f2sdram~O_BONDING_OUT_10 ;
wire \f2sdram~O_BONDING_OUT_11 ;
wire \f2sdram~O_BONDING_OUT_12 ;
wire \f2sdram~O_BONDING_OUT_13 ;
wire \clocks_resets~h2f_cold_rst_n ;
wire \h2f_ARADDR[9] ;
wire \h2f_ARADDR[10] ;
wire \h2f_ARADDR[11] ;
wire \h2f_ARADDR[12] ;
wire \h2f_ARADDR[13] ;
wire \h2f_ARADDR[14] ;
wire \h2f_ARADDR[15] ;
wire \h2f_ARADDR[16] ;
wire \h2f_ARADDR[17] ;
wire \h2f_ARADDR[18] ;
wire \h2f_ARADDR[19] ;
wire \h2f_ARADDR[20] ;
wire \h2f_ARADDR[21] ;
wire \h2f_ARADDR[22] ;
wire \h2f_ARADDR[23] ;
wire \h2f_ARADDR[24] ;
wire \h2f_ARADDR[25] ;
wire \h2f_ARADDR[26] ;
wire \h2f_ARADDR[27] ;
wire \h2f_ARADDR[28] ;
wire \h2f_ARADDR[29] ;

wire [31:0] tpiu_TRACE_DATA_bus;
wire [3:0] f2sdram_BONDING_OUT_1_bus;
wire [29:0] hps2fpga_ARADDR_bus;
wire [1:0] hps2fpga_ARBURST_bus;
wire [11:0] hps2fpga_ARID_bus;
wire [3:0] hps2fpga_ARLEN_bus;
wire [2:0] hps2fpga_ARSIZE_bus;
wire [29:0] hps2fpga_AWADDR_bus;
wire [1:0] hps2fpga_AWBURST_bus;
wire [11:0] hps2fpga_AWID_bus;
wire [3:0] hps2fpga_AWLEN_bus;
wire [2:0] hps2fpga_AWSIZE_bus;
wire [127:0] hps2fpga_WDATA_bus;
wire [15:0] hps2fpga_WSTRB_bus;

assign \tpiu~trace_data  = tpiu_TRACE_DATA_bus[0];
assign \tpiu~O_TRACE_DATA1  = tpiu_TRACE_DATA_bus[1];
assign \tpiu~O_TRACE_DATA2  = tpiu_TRACE_DATA_bus[2];
assign \tpiu~O_TRACE_DATA3  = tpiu_TRACE_DATA_bus[3];
assign \tpiu~O_TRACE_DATA4  = tpiu_TRACE_DATA_bus[4];
assign \tpiu~O_TRACE_DATA5  = tpiu_TRACE_DATA_bus[5];
assign \tpiu~O_TRACE_DATA6  = tpiu_TRACE_DATA_bus[6];
assign \tpiu~O_TRACE_DATA7  = tpiu_TRACE_DATA_bus[7];
assign \tpiu~O_TRACE_DATA8  = tpiu_TRACE_DATA_bus[8];
assign \tpiu~O_TRACE_DATA9  = tpiu_TRACE_DATA_bus[9];
assign \tpiu~O_TRACE_DATA10  = tpiu_TRACE_DATA_bus[10];
assign \tpiu~O_TRACE_DATA11  = tpiu_TRACE_DATA_bus[11];
assign \tpiu~O_TRACE_DATA12  = tpiu_TRACE_DATA_bus[12];
assign \tpiu~O_TRACE_DATA13  = tpiu_TRACE_DATA_bus[13];
assign \tpiu~O_TRACE_DATA14  = tpiu_TRACE_DATA_bus[14];
assign \tpiu~O_TRACE_DATA15  = tpiu_TRACE_DATA_bus[15];
assign \tpiu~O_TRACE_DATA16  = tpiu_TRACE_DATA_bus[16];
assign \tpiu~O_TRACE_DATA17  = tpiu_TRACE_DATA_bus[17];
assign \tpiu~O_TRACE_DATA18  = tpiu_TRACE_DATA_bus[18];
assign \tpiu~O_TRACE_DATA19  = tpiu_TRACE_DATA_bus[19];
assign \tpiu~O_TRACE_DATA20  = tpiu_TRACE_DATA_bus[20];
assign \tpiu~O_TRACE_DATA21  = tpiu_TRACE_DATA_bus[21];
assign \tpiu~O_TRACE_DATA22  = tpiu_TRACE_DATA_bus[22];
assign \tpiu~O_TRACE_DATA23  = tpiu_TRACE_DATA_bus[23];
assign \tpiu~O_TRACE_DATA24  = tpiu_TRACE_DATA_bus[24];
assign \tpiu~O_TRACE_DATA25  = tpiu_TRACE_DATA_bus[25];
assign \tpiu~O_TRACE_DATA26  = tpiu_TRACE_DATA_bus[26];
assign \tpiu~O_TRACE_DATA27  = tpiu_TRACE_DATA_bus[27];
assign \tpiu~O_TRACE_DATA28  = tpiu_TRACE_DATA_bus[28];
assign \tpiu~O_TRACE_DATA29  = tpiu_TRACE_DATA_bus[29];
assign \tpiu~O_TRACE_DATA30  = tpiu_TRACE_DATA_bus[30];
assign \tpiu~O_TRACE_DATA31  = tpiu_TRACE_DATA_bus[31];

assign \f2sdram~O_BONDING_OUT_10  = f2sdram_BONDING_OUT_1_bus[0];
assign \f2sdram~O_BONDING_OUT_11  = f2sdram_BONDING_OUT_1_bus[1];
assign \f2sdram~O_BONDING_OUT_12  = f2sdram_BONDING_OUT_1_bus[2];
assign \f2sdram~O_BONDING_OUT_13  = f2sdram_BONDING_OUT_1_bus[3];

assign h2f_ARADDR[0] = hps2fpga_ARADDR_bus[0];
assign h2f_ARADDR[1] = hps2fpga_ARADDR_bus[1];
assign h2f_ARADDR[2] = hps2fpga_ARADDR_bus[2];
assign h2f_ARADDR[3] = hps2fpga_ARADDR_bus[3];
assign h2f_ARADDR[4] = hps2fpga_ARADDR_bus[4];
assign h2f_ARADDR[5] = hps2fpga_ARADDR_bus[5];
assign h2f_ARADDR[6] = hps2fpga_ARADDR_bus[6];
assign h2f_ARADDR[7] = hps2fpga_ARADDR_bus[7];
assign h2f_ARADDR[8] = hps2fpga_ARADDR_bus[8];
assign \h2f_ARADDR[9]  = hps2fpga_ARADDR_bus[9];
assign \h2f_ARADDR[10]  = hps2fpga_ARADDR_bus[10];
assign \h2f_ARADDR[11]  = hps2fpga_ARADDR_bus[11];
assign \h2f_ARADDR[12]  = hps2fpga_ARADDR_bus[12];
assign \h2f_ARADDR[13]  = hps2fpga_ARADDR_bus[13];
assign \h2f_ARADDR[14]  = hps2fpga_ARADDR_bus[14];
assign \h2f_ARADDR[15]  = hps2fpga_ARADDR_bus[15];
assign \h2f_ARADDR[16]  = hps2fpga_ARADDR_bus[16];
assign \h2f_ARADDR[17]  = hps2fpga_ARADDR_bus[17];
assign \h2f_ARADDR[18]  = hps2fpga_ARADDR_bus[18];
assign \h2f_ARADDR[19]  = hps2fpga_ARADDR_bus[19];
assign \h2f_ARADDR[20]  = hps2fpga_ARADDR_bus[20];
assign \h2f_ARADDR[21]  = hps2fpga_ARADDR_bus[21];
assign \h2f_ARADDR[22]  = hps2fpga_ARADDR_bus[22];
assign \h2f_ARADDR[23]  = hps2fpga_ARADDR_bus[23];
assign \h2f_ARADDR[24]  = hps2fpga_ARADDR_bus[24];
assign \h2f_ARADDR[25]  = hps2fpga_ARADDR_bus[25];
assign \h2f_ARADDR[26]  = hps2fpga_ARADDR_bus[26];
assign \h2f_ARADDR[27]  = hps2fpga_ARADDR_bus[27];
assign \h2f_ARADDR[28]  = hps2fpga_ARADDR_bus[28];
assign \h2f_ARADDR[29]  = hps2fpga_ARADDR_bus[29];

assign h2f_ARBURST[0] = hps2fpga_ARBURST_bus[0];
assign h2f_ARBURST[1] = hps2fpga_ARBURST_bus[1];

assign h2f_ARID[0] = hps2fpga_ARID_bus[0];
assign h2f_ARID[1] = hps2fpga_ARID_bus[1];
assign h2f_ARID[2] = hps2fpga_ARID_bus[2];
assign h2f_ARID[3] = hps2fpga_ARID_bus[3];
assign h2f_ARID[4] = hps2fpga_ARID_bus[4];
assign h2f_ARID[5] = hps2fpga_ARID_bus[5];
assign h2f_ARID[6] = hps2fpga_ARID_bus[6];
assign h2f_ARID[7] = hps2fpga_ARID_bus[7];
assign h2f_ARID[8] = hps2fpga_ARID_bus[8];
assign h2f_ARID[9] = hps2fpga_ARID_bus[9];
assign h2f_ARID[10] = hps2fpga_ARID_bus[10];
assign h2f_ARID[11] = hps2fpga_ARID_bus[11];

assign h2f_ARLEN[0] = hps2fpga_ARLEN_bus[0];
assign h2f_ARLEN[1] = hps2fpga_ARLEN_bus[1];
assign h2f_ARLEN[2] = hps2fpga_ARLEN_bus[2];
assign h2f_ARLEN[3] = hps2fpga_ARLEN_bus[3];

assign h2f_ARSIZE[0] = hps2fpga_ARSIZE_bus[0];
assign h2f_ARSIZE[1] = hps2fpga_ARSIZE_bus[1];
assign h2f_ARSIZE[2] = hps2fpga_ARSIZE_bus[2];

assign h2f_AWADDR[0] = hps2fpga_AWADDR_bus[0];
assign h2f_AWADDR[1] = hps2fpga_AWADDR_bus[1];
assign h2f_AWADDR[2] = hps2fpga_AWADDR_bus[2];
assign h2f_AWADDR[3] = hps2fpga_AWADDR_bus[3];
assign h2f_AWADDR[4] = hps2fpga_AWADDR_bus[4];
assign h2f_AWADDR[5] = hps2fpga_AWADDR_bus[5];
assign h2f_AWADDR[6] = hps2fpga_AWADDR_bus[6];
assign h2f_AWADDR[7] = hps2fpga_AWADDR_bus[7];
assign h2f_AWADDR[8] = hps2fpga_AWADDR_bus[8];

assign h2f_AWBURST[0] = hps2fpga_AWBURST_bus[0];
assign h2f_AWBURST[1] = hps2fpga_AWBURST_bus[1];

assign h2f_AWID[0] = hps2fpga_AWID_bus[0];
assign h2f_AWID[1] = hps2fpga_AWID_bus[1];
assign h2f_AWID[2] = hps2fpga_AWID_bus[2];
assign h2f_AWID[3] = hps2fpga_AWID_bus[3];
assign h2f_AWID[4] = hps2fpga_AWID_bus[4];
assign h2f_AWID[5] = hps2fpga_AWID_bus[5];
assign h2f_AWID[6] = hps2fpga_AWID_bus[6];
assign h2f_AWID[7] = hps2fpga_AWID_bus[7];
assign h2f_AWID[8] = hps2fpga_AWID_bus[8];
assign h2f_AWID[9] = hps2fpga_AWID_bus[9];
assign h2f_AWID[10] = hps2fpga_AWID_bus[10];
assign h2f_AWID[11] = hps2fpga_AWID_bus[11];

assign h2f_AWLEN[0] = hps2fpga_AWLEN_bus[0];
assign h2f_AWLEN[1] = hps2fpga_AWLEN_bus[1];
assign h2f_AWLEN[2] = hps2fpga_AWLEN_bus[2];
assign h2f_AWLEN[3] = hps2fpga_AWLEN_bus[3];

assign h2f_AWSIZE[0] = hps2fpga_AWSIZE_bus[0];
assign h2f_AWSIZE[1] = hps2fpga_AWSIZE_bus[1];
assign h2f_AWSIZE[2] = hps2fpga_AWSIZE_bus[2];

assign h2f_WDATA[0] = hps2fpga_WDATA_bus[0];
assign h2f_WDATA[1] = hps2fpga_WDATA_bus[1];
assign h2f_WDATA[2] = hps2fpga_WDATA_bus[2];
assign h2f_WDATA[3] = hps2fpga_WDATA_bus[3];
assign h2f_WDATA[4] = hps2fpga_WDATA_bus[4];
assign h2f_WDATA[5] = hps2fpga_WDATA_bus[5];
assign h2f_WDATA[6] = hps2fpga_WDATA_bus[6];
assign h2f_WDATA[7] = hps2fpga_WDATA_bus[7];
assign h2f_WDATA[8] = hps2fpga_WDATA_bus[8];

assign h2f_WSTRB[0] = hps2fpga_WSTRB_bus[0];
assign h2f_WSTRB[1] = hps2fpga_WSTRB_bus[1];
assign h2f_WSTRB[2] = hps2fpga_WSTRB_bus[2];
assign h2f_WSTRB[3] = hps2fpga_WSTRB_bus[3];

cyclonev_hps_interface_clocks_resets clocks_resets(
	.f2h_cold_rst_req_n(vcc),
	.f2h_dbg_rst_req_n(vcc),
	.f2h_pending_rst_ack(vcc),
	.f2h_periph_ref_clk(gnd),
	.f2h_sdram_ref_clk(gnd),
	.f2h_warm_rst_req_n(vcc),
	.ptp_ref_clk(gnd),
	.h2f_cold_rst_n(\clocks_resets~h2f_cold_rst_n ),
	.h2f_pending_rst_req_n(),
	.h2f_rst_n(h2f_rst_n[0]),
	.h2f_user0_clk(),
	.h2f_user1_clk(),
	.h2f_user2_clk());
defparam clocks_resets.h2f_user0_clk_freq = 100;
defparam clocks_resets.h2f_user1_clk_freq = 100;
defparam clocks_resets.h2f_user2_clk_freq = 100;

cyclonev_hps_interface_hps2fpga hps2fpga(
	.arready(h2f_ARREADY[0]),
	.awready(h2f_AWREADY[0]),
	.bvalid(h2f_BVALID[0]),
	.clk(h2f_axi_clk[0]),
	.rlast(h2f_RLAST[0]),
	.rvalid(h2f_RVALID[0]),
	.wready(h2f_WREADY[0]),
	.bid({h2f_BID[11],h2f_BID[10],h2f_BID[9],h2f_BID[8],h2f_BID[7],h2f_BID[6],h2f_BID[5],h2f_BID[4],h2f_BID[3],h2f_BID[2],h2f_BID[1],h2f_BID[0]}),
	.bresp({gnd,gnd}),
	.port_size_config({gnd,gnd}),
	.rdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,h2f_RDATA[10],h2f_RDATA[9],h2f_RDATA[8],h2f_RDATA[7],h2f_RDATA[6],h2f_RDATA[5],h2f_RDATA[4],h2f_RDATA[3],h2f_RDATA[2],h2f_RDATA[1],h2f_RDATA[0]}),
	.rid({h2f_RID[11],h2f_RID[10],h2f_RID[9],h2f_RID[8],h2f_RID[7],h2f_RID[6],h2f_RID[5],h2f_RID[4],h2f_RID[3],h2f_RID[2],h2f_RID[1],h2f_RID[0]}),
	.rresp({gnd,gnd}),
	.arvalid(h2f_ARVALID[0]),
	.awvalid(h2f_AWVALID[0]),
	.bready(h2f_BREADY[0]),
	.rready(h2f_RREADY[0]),
	.wlast(h2f_WLAST[0]),
	.wvalid(h2f_WVALID[0]),
	.araddr(hps2fpga_ARADDR_bus),
	.arburst(hps2fpga_ARBURST_bus),
	.arcache(),
	.arid(hps2fpga_ARID_bus),
	.arlen(hps2fpga_ARLEN_bus),
	.arlock(),
	.arprot(),
	.arsize(hps2fpga_ARSIZE_bus),
	.awaddr(hps2fpga_AWADDR_bus),
	.awburst(hps2fpga_AWBURST_bus),
	.awcache(),
	.awid(hps2fpga_AWID_bus),
	.awlen(hps2fpga_AWLEN_bus),
	.awlock(),
	.awprot(),
	.awsize(hps2fpga_AWSIZE_bus),
	.wdata(hps2fpga_WDATA_bus),
	.wid(),
	.wstrb(hps2fpga_WSTRB_bus));
defparam hps2fpga.data_width = 32;

cyclonev_hps_interface_dbg_apb debug_apb(
	.p_slv_err(gnd),
	.p_ready(gnd),
	.p_clk(gnd),
	.p_clk_en(gnd),
	.dbg_apb_disable(gnd),
	.p_rdata(32'b00000000000000000000000000000000),
	.p_addr_31(\debug_apb~O_P_ADDR_31 ),
	.p_write(),
	.p_sel(),
	.p_enable(),
	.p_reset_n(),
	.p_addr(),
	.p_wdata());
defparam debug_apb.dummy_param = 256;

cyclonev_hps_interface_tpiu_trace tpiu(
	.traceclk_ctl(vcc),
	.traceclkin(gnd),
	.traceclk(),
	.trace_data(tpiu_TRACE_DATA_bus));

cyclonev_hps_interface_boot_from_fpga boot_from_fpga(
	.boot_from_fpga_on_failure(gnd),
	.boot_from_fpga_ready(gnd),
	.bsel_en(gnd),
	.csel_en(gnd),
	.bsel({gnd,gnd,vcc}),
	.csel({gnd,vcc}),
	.fake_dout(\boot_from_fpga~fake_dout ));

cyclonev_hps_interface_fpga2hps fpga2hps(
	.arvalid(gnd),
	.awvalid(gnd),
	.bready(gnd),
	.clk(gnd),
	.rready(gnd),
	.wlast(gnd),
	.wvalid(gnd),
	.araddr(32'b00000000000000000000000000000000),
	.arburst(2'b00),
	.arcache(4'b0000),
	.arid(8'b00000000),
	.arlen(4'b0000),
	.arlock(2'b00),
	.arprot(3'b000),
	.arsize(3'b000),
	.aruser(5'b00000),
	.awaddr(32'b00000000000000000000000000000000),
	.awburst(2'b00),
	.awcache(4'b0000),
	.awid(8'b00000000),
	.awlen(4'b0000),
	.awlock(2'b00),
	.awprot(3'b000),
	.awsize(3'b000),
	.awuser(5'b00000),
	.port_size_config({vcc,vcc}),
	.wdata(128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
	.wid(8'b00000000),
	.wstrb(16'b0000000000000000),
	.arready(\fpga2hps~arready ),
	.awready(),
	.bvalid(),
	.rlast(),
	.rvalid(),
	.wready(),
	.bid(),
	.bresp(),
	.rdata(),
	.rid(),
	.rresp());
defparam fpga2hps.data_width = 32;

cyclonev_hps_interface_fpga2sdram f2sdram(
	.cmd_port_clk_0(gnd),
	.cmd_port_clk_1(gnd),
	.cmd_port_clk_2(gnd),
	.cmd_port_clk_3(gnd),
	.cmd_port_clk_4(gnd),
	.cmd_port_clk_5(gnd),
	.cmd_valid_0(gnd),
	.cmd_valid_1(gnd),
	.cmd_valid_2(gnd),
	.cmd_valid_3(gnd),
	.cmd_valid_4(gnd),
	.cmd_valid_5(gnd),
	.rd_clk_0(gnd),
	.rd_clk_1(gnd),
	.rd_clk_2(gnd),
	.rd_clk_3(gnd),
	.rd_ready_0(gnd),
	.rd_ready_1(gnd),
	.rd_ready_2(gnd),
	.rd_ready_3(gnd),
	.wr_clk_0(gnd),
	.wr_clk_1(gnd),
	.wr_clk_2(gnd),
	.wr_clk_3(gnd),
	.wr_valid_0(gnd),
	.wr_valid_1(gnd),
	.wr_valid_2(gnd),
	.wr_valid_3(gnd),
	.wrack_ready_0(gnd),
	.wrack_ready_1(gnd),
	.wrack_ready_2(gnd),
	.wrack_ready_3(gnd),
	.wrack_ready_4(gnd),
	.wrack_ready_5(gnd),
	.cfg_axi_mm_select({gnd,gnd,gnd,gnd,gnd,gnd}),
	.cfg_cport_rfifo_map({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.cfg_cport_type({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.cfg_cport_wfifo_map({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.cfg_port_width({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.cfg_rfifo_cport_map({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.cfg_wfifo_cport_map({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.cmd_data_0(60'b000000000000000000000000000000000000000000000000000000000000),
	.cmd_data_1(60'b000000000000000000000000000000000000000000000000000000000000),
	.cmd_data_2(60'b000000000000000000000000000000000000000000000000000000000000),
	.cmd_data_3(60'b000000000000000000000000000000000000000000000000000000000000),
	.cmd_data_4(60'b000000000000000000000000000000000000000000000000000000000000),
	.cmd_data_5(60'b000000000000000000000000000000000000000000000000000000000000),
	.wr_data_0(90'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
	.wr_data_1(90'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
	.wr_data_2(90'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
	.wr_data_3(90'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
	.cmd_ready_0(),
	.cmd_ready_1(),
	.cmd_ready_2(),
	.cmd_ready_3(),
	.cmd_ready_4(),
	.cmd_ready_5(),
	.rd_valid_0(),
	.rd_valid_1(),
	.rd_valid_2(),
	.rd_valid_3(),
	.wr_ready_0(),
	.wr_ready_1(),
	.wr_ready_2(),
	.wr_ready_3(),
	.wrack_valid_0(),
	.wrack_valid_1(),
	.wrack_valid_2(),
	.wrack_valid_3(),
	.wrack_valid_4(),
	.wrack_valid_5(),
	.bonding_out_1(f2sdram_BONDING_OUT_1_bus),
	.bonding_out_2(),
	.rd_data_0(),
	.rd_data_1(),
	.rd_data_2(),
	.rd_data_3(),
	.wrack_data_0(),
	.wrack_data_1(),
	.wrack_data_2(),
	.wrack_data_3(),
	.wrack_data_4(),
	.wrack_data_5());

endmodule

module spw_babasu_spw_babasu_mm_interconnect_0 (
	h2f_ARVALID_0,
	h2f_AWVALID_0,
	h2f_BREADY_0,
	h2f_RREADY_0,
	h2f_WLAST_0,
	h2f_WVALID_0,
	h2f_ARADDR_0,
	h2f_ARADDR_1,
	h2f_ARADDR_2,
	h2f_ARADDR_3,
	h2f_ARADDR_4,
	h2f_ARADDR_5,
	h2f_ARADDR_6,
	h2f_ARADDR_7,
	h2f_ARADDR_8,
	h2f_ARBURST_0,
	h2f_ARBURST_1,
	h2f_ARID_0,
	h2f_ARID_1,
	h2f_ARID_2,
	h2f_ARID_3,
	h2f_ARID_4,
	h2f_ARID_5,
	h2f_ARID_6,
	h2f_ARID_7,
	h2f_ARID_8,
	h2f_ARID_9,
	h2f_ARID_10,
	h2f_ARID_11,
	h2f_ARLEN_0,
	h2f_ARLEN_1,
	h2f_ARLEN_2,
	h2f_ARLEN_3,
	h2f_ARSIZE_0,
	h2f_ARSIZE_1,
	h2f_ARSIZE_2,
	h2f_AWADDR_0,
	h2f_AWADDR_1,
	h2f_AWADDR_2,
	h2f_AWADDR_3,
	h2f_AWADDR_4,
	h2f_AWADDR_5,
	h2f_AWADDR_6,
	h2f_AWADDR_7,
	h2f_AWADDR_8,
	h2f_AWBURST_0,
	h2f_AWBURST_1,
	h2f_AWID_0,
	h2f_AWID_1,
	h2f_AWID_2,
	h2f_AWID_3,
	h2f_AWID_4,
	h2f_AWID_5,
	h2f_AWID_6,
	h2f_AWID_7,
	h2f_AWID_8,
	h2f_AWID_9,
	h2f_AWID_10,
	h2f_AWID_11,
	h2f_AWLEN_0,
	h2f_AWLEN_1,
	h2f_AWLEN_2,
	h2f_AWLEN_3,
	h2f_AWSIZE_0,
	h2f_AWSIZE_1,
	h2f_AWSIZE_2,
	h2f_WDATA_0,
	h2f_WDATA_1,
	h2f_WDATA_2,
	h2f_WDATA_3,
	h2f_WDATA_4,
	h2f_WDATA_5,
	h2f_WDATA_6,
	h2f_WDATA_7,
	h2f_WDATA_8,
	h2f_WSTRB_0,
	h2f_WSTRB_1,
	h2f_WSTRB_2,
	h2f_WSTRB_3,
	wait_latency_counter_1,
	wait_latency_counter_0,
	wait_latency_counter_11,
	wait_latency_counter_01,
	wait_latency_counter_12,
	wait_latency_counter_02,
	wait_latency_counter_13,
	wait_latency_counter_03,
	wait_latency_counter_14,
	wait_latency_counter_04,
	wait_latency_counter_15,
	wait_latency_counter_05,
	wait_latency_counter_16,
	wait_latency_counter_06,
	wait_latency_counter_17,
	wait_latency_counter_07,
	wait_latency_counter_18,
	wait_latency_counter_08,
	wait_latency_counter_19,
	wait_latency_counter_09,
	cmd_sink_ready,
	nonposted_cmd_accepted,
	WideOr1,
	src_payload_0,
	WideOr11,
	nonposted_cmd_accepted1,
	src_data_105,
	src_data_106,
	src_data_107,
	src_data_108,
	src_data_109,
	src_data_110,
	src_data_111,
	src_data_112,
	src_data_113,
	src_data_114,
	src_data_115,
	src_data_116,
	src_data_0,
	src_payload,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_data_1051,
	src_data_1061,
	src_data_1071,
	src_data_1081,
	src_data_1091,
	src_data_1101,
	src_data_1111,
	src_data_1121,
	src_data_1131,
	src_data_1141,
	src_data_1151,
	src_data_1161,
	m0_write,
	in_data_reg_0,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	altera_reset_synchronizer_int_chain_out,
	in_data_reg_01,
	m0_write1,
	int_nxt_addr_reg_dly_31,
	int_nxt_addr_reg_dly_21,
	in_data_reg_1,
	in_data_reg_2,
	in_data_reg_3,
	in_data_reg_4,
	in_data_reg_5,
	in_data_reg_6,
	in_data_reg_7,
	in_data_reg_8,
	m0_write2,
	in_data_reg_02,
	int_nxt_addr_reg_dly_32,
	int_nxt_addr_reg_dly_22,
	m0_write3,
	in_data_reg_03,
	int_nxt_addr_reg_dly_33,
	int_nxt_addr_reg_dly_23,
	m0_write4,
	in_data_reg_04,
	int_nxt_addr_reg_dly_34,
	int_nxt_addr_reg_dly_24,
	m0_write5,
	in_data_reg_05,
	int_nxt_addr_reg_dly_35,
	int_nxt_addr_reg_dly_25,
	m0_write6,
	in_data_reg_06,
	int_nxt_addr_reg_dly_36,
	int_nxt_addr_reg_dly_26,
	in_data_reg_07,
	m0_write7,
	int_nxt_addr_reg_dly_37,
	int_nxt_addr_reg_dly_27,
	in_data_reg_11,
	in_data_reg_21,
	in_data_reg_31,
	in_data_reg_41,
	in_data_reg_51,
	in_data_reg_61,
	in_data_reg_71,
	in_data_reg_08,
	m0_write8,
	int_nxt_addr_reg_dly_38,
	int_nxt_addr_reg_dly_28,
	in_data_reg_12,
	in_data_reg_22,
	in_data_reg_32,
	in_data_reg_42,
	in_data_reg_52,
	in_data_reg_62,
	m0_write9,
	in_data_reg_09,
	int_nxt_addr_reg_dly_39,
	int_nxt_addr_reg_dly_29,
	altera_reset_synchronizer_int_chain_out1,
	readdata_0,
	readdata_01,
	readdata_02,
	readdata_03,
	readdata_04,
	readdata_05,
	readdata_06,
	readdata_07,
	readdata_08,
	readdata_09,
	readdata_010,
	readdata_011,
	readdata_012,
	readdata_013,
	readdata_014,
	readdata_015,
	readdata_016,
	readdata_1,
	readdata_11,
	readdata_12,
	readdata_13,
	readdata_14,
	readdata_15,
	readdata_16,
	readdata_2,
	readdata_21,
	readdata_22,
	readdata_23,
	readdata_24,
	readdata_25,
	readdata_26,
	readdata_3,
	readdata_31,
	readdata_32,
	readdata_33,
	readdata_34,
	readdata_35,
	readdata_4,
	readdata_41,
	readdata_42,
	readdata_43,
	readdata_44,
	readdata_45,
	readdata_5,
	readdata_51,
	readdata_52,
	readdata_53,
	readdata_54,
	readdata_55,
	readdata_6,
	readdata_61,
	readdata_62,
	readdata_63,
	readdata_64,
	readdata_65,
	readdata_7,
	readdata_71,
	readdata_72,
	readdata_73,
	readdata_74,
	readdata_8,
	readdata_81,
	readdata_82,
	readdata_9,
	readdata_10,
	int_nxt_addr_reg_dly_310,
	int_nxt_addr_reg_dly_210,
	int_nxt_addr_reg_dly_311,
	int_nxt_addr_reg_dly_211,
	int_nxt_addr_reg_dly_312,
	int_nxt_addr_reg_dly_212,
	int_nxt_addr_reg_dly_313,
	int_nxt_addr_reg_dly_213,
	int_nxt_addr_reg_dly_314,
	int_nxt_addr_reg_dly_214,
	int_nxt_addr_reg_dly_315,
	int_nxt_addr_reg_dly_215,
	int_nxt_addr_reg_dly_316,
	int_nxt_addr_reg_dly_216,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARVALID_0;
input 	h2f_AWVALID_0;
input 	h2f_BREADY_0;
input 	h2f_RREADY_0;
input 	h2f_WLAST_0;
input 	h2f_WVALID_0;
input 	h2f_ARADDR_0;
input 	h2f_ARADDR_1;
input 	h2f_ARADDR_2;
input 	h2f_ARADDR_3;
input 	h2f_ARADDR_4;
input 	h2f_ARADDR_5;
input 	h2f_ARADDR_6;
input 	h2f_ARADDR_7;
input 	h2f_ARADDR_8;
input 	h2f_ARBURST_0;
input 	h2f_ARBURST_1;
input 	h2f_ARID_0;
input 	h2f_ARID_1;
input 	h2f_ARID_2;
input 	h2f_ARID_3;
input 	h2f_ARID_4;
input 	h2f_ARID_5;
input 	h2f_ARID_6;
input 	h2f_ARID_7;
input 	h2f_ARID_8;
input 	h2f_ARID_9;
input 	h2f_ARID_10;
input 	h2f_ARID_11;
input 	h2f_ARLEN_0;
input 	h2f_ARLEN_1;
input 	h2f_ARLEN_2;
input 	h2f_ARLEN_3;
input 	h2f_ARSIZE_0;
input 	h2f_ARSIZE_1;
input 	h2f_ARSIZE_2;
input 	h2f_AWADDR_0;
input 	h2f_AWADDR_1;
input 	h2f_AWADDR_2;
input 	h2f_AWADDR_3;
input 	h2f_AWADDR_4;
input 	h2f_AWADDR_5;
input 	h2f_AWADDR_6;
input 	h2f_AWADDR_7;
input 	h2f_AWADDR_8;
input 	h2f_AWBURST_0;
input 	h2f_AWBURST_1;
input 	h2f_AWID_0;
input 	h2f_AWID_1;
input 	h2f_AWID_2;
input 	h2f_AWID_3;
input 	h2f_AWID_4;
input 	h2f_AWID_5;
input 	h2f_AWID_6;
input 	h2f_AWID_7;
input 	h2f_AWID_8;
input 	h2f_AWID_9;
input 	h2f_AWID_10;
input 	h2f_AWID_11;
input 	h2f_AWLEN_0;
input 	h2f_AWLEN_1;
input 	h2f_AWLEN_2;
input 	h2f_AWLEN_3;
input 	h2f_AWSIZE_0;
input 	h2f_AWSIZE_1;
input 	h2f_AWSIZE_2;
input 	h2f_WDATA_0;
input 	h2f_WDATA_1;
input 	h2f_WDATA_2;
input 	h2f_WDATA_3;
input 	h2f_WDATA_4;
input 	h2f_WDATA_5;
input 	h2f_WDATA_6;
input 	h2f_WDATA_7;
input 	h2f_WDATA_8;
input 	h2f_WSTRB_0;
input 	h2f_WSTRB_1;
input 	h2f_WSTRB_2;
input 	h2f_WSTRB_3;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
output 	wait_latency_counter_11;
output 	wait_latency_counter_01;
output 	wait_latency_counter_12;
output 	wait_latency_counter_02;
output 	wait_latency_counter_13;
output 	wait_latency_counter_03;
output 	wait_latency_counter_14;
output 	wait_latency_counter_04;
output 	wait_latency_counter_15;
output 	wait_latency_counter_05;
output 	wait_latency_counter_16;
output 	wait_latency_counter_06;
output 	wait_latency_counter_17;
output 	wait_latency_counter_07;
output 	wait_latency_counter_18;
output 	wait_latency_counter_08;
output 	wait_latency_counter_19;
output 	wait_latency_counter_09;
output 	cmd_sink_ready;
output 	nonposted_cmd_accepted;
output 	WideOr1;
output 	src_payload_0;
output 	WideOr11;
output 	nonposted_cmd_accepted1;
output 	src_data_105;
output 	src_data_106;
output 	src_data_107;
output 	src_data_108;
output 	src_data_109;
output 	src_data_110;
output 	src_data_111;
output 	src_data_112;
output 	src_data_113;
output 	src_data_114;
output 	src_data_115;
output 	src_data_116;
output 	src_data_0;
output 	src_payload;
output 	src_payload1;
output 	src_payload2;
output 	src_payload3;
output 	src_payload4;
output 	src_payload5;
output 	src_payload6;
output 	src_payload7;
output 	src_payload8;
output 	src_payload9;
output 	src_data_1051;
output 	src_data_1061;
output 	src_data_1071;
output 	src_data_1081;
output 	src_data_1091;
output 	src_data_1101;
output 	src_data_1111;
output 	src_data_1121;
output 	src_data_1131;
output 	src_data_1141;
output 	src_data_1151;
output 	src_data_1161;
output 	m0_write;
output 	in_data_reg_0;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
input 	altera_reset_synchronizer_int_chain_out;
output 	in_data_reg_01;
output 	m0_write1;
output 	int_nxt_addr_reg_dly_31;
output 	int_nxt_addr_reg_dly_21;
output 	in_data_reg_1;
output 	in_data_reg_2;
output 	in_data_reg_3;
output 	in_data_reg_4;
output 	in_data_reg_5;
output 	in_data_reg_6;
output 	in_data_reg_7;
output 	in_data_reg_8;
output 	m0_write2;
output 	in_data_reg_02;
output 	int_nxt_addr_reg_dly_32;
output 	int_nxt_addr_reg_dly_22;
output 	m0_write3;
output 	in_data_reg_03;
output 	int_nxt_addr_reg_dly_33;
output 	int_nxt_addr_reg_dly_23;
output 	m0_write4;
output 	in_data_reg_04;
output 	int_nxt_addr_reg_dly_34;
output 	int_nxt_addr_reg_dly_24;
output 	m0_write5;
output 	in_data_reg_05;
output 	int_nxt_addr_reg_dly_35;
output 	int_nxt_addr_reg_dly_25;
output 	m0_write6;
output 	in_data_reg_06;
output 	int_nxt_addr_reg_dly_36;
output 	int_nxt_addr_reg_dly_26;
output 	in_data_reg_07;
output 	m0_write7;
output 	int_nxt_addr_reg_dly_37;
output 	int_nxt_addr_reg_dly_27;
output 	in_data_reg_11;
output 	in_data_reg_21;
output 	in_data_reg_31;
output 	in_data_reg_41;
output 	in_data_reg_51;
output 	in_data_reg_61;
output 	in_data_reg_71;
output 	in_data_reg_08;
output 	m0_write8;
output 	int_nxt_addr_reg_dly_38;
output 	int_nxt_addr_reg_dly_28;
output 	in_data_reg_12;
output 	in_data_reg_22;
output 	in_data_reg_32;
output 	in_data_reg_42;
output 	in_data_reg_52;
output 	in_data_reg_62;
output 	m0_write9;
output 	in_data_reg_09;
output 	int_nxt_addr_reg_dly_39;
output 	int_nxt_addr_reg_dly_29;
input 	altera_reset_synchronizer_int_chain_out1;
input 	readdata_0;
input 	readdata_01;
input 	readdata_02;
input 	readdata_03;
input 	readdata_04;
input 	readdata_05;
input 	readdata_06;
input 	readdata_07;
input 	readdata_08;
input 	readdata_09;
input 	readdata_010;
input 	readdata_011;
input 	readdata_012;
input 	readdata_013;
input 	readdata_014;
input 	readdata_015;
input 	readdata_016;
input 	readdata_1;
input 	readdata_11;
input 	readdata_12;
input 	readdata_13;
input 	readdata_14;
input 	readdata_15;
input 	readdata_16;
input 	readdata_2;
input 	readdata_21;
input 	readdata_22;
input 	readdata_23;
input 	readdata_24;
input 	readdata_25;
input 	readdata_26;
input 	readdata_3;
input 	readdata_31;
input 	readdata_32;
input 	readdata_33;
input 	readdata_34;
input 	readdata_35;
input 	readdata_4;
input 	readdata_41;
input 	readdata_42;
input 	readdata_43;
input 	readdata_44;
input 	readdata_45;
input 	readdata_5;
input 	readdata_51;
input 	readdata_52;
input 	readdata_53;
input 	readdata_54;
input 	readdata_55;
input 	readdata_6;
input 	readdata_61;
input 	readdata_62;
input 	readdata_63;
input 	readdata_64;
input 	readdata_65;
input 	readdata_7;
input 	readdata_71;
input 	readdata_72;
input 	readdata_73;
input 	readdata_74;
input 	readdata_8;
input 	readdata_81;
input 	readdata_82;
input 	readdata_9;
input 	readdata_10;
output 	int_nxt_addr_reg_dly_310;
output 	int_nxt_addr_reg_dly_210;
output 	int_nxt_addr_reg_dly_311;
output 	int_nxt_addr_reg_dly_211;
output 	int_nxt_addr_reg_dly_312;
output 	int_nxt_addr_reg_dly_212;
output 	int_nxt_addr_reg_dly_313;
output 	int_nxt_addr_reg_dly_213;
output 	int_nxt_addr_reg_dly_314;
output 	int_nxt_addr_reg_dly_214;
output 	int_nxt_addr_reg_dly_315;
output 	int_nxt_addr_reg_dly_215;
output 	int_nxt_addr_reg_dly_316;
output 	int_nxt_addr_reg_dly_216;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \hps_0_h2f_axi_master_agent|align_address_to_size|address_burst[8]~q ;
wire \hps_0_h2f_axi_master_agent|align_address_to_size|address_burst[7]~q ;
wire \hps_0_h2f_axi_master_agent|align_address_to_size|address_burst[6]~q ;
wire \hps_0_h2f_axi_master_agent|Add5~1_sumout ;
wire \hps_0_h2f_axi_master_agent|Add5~5_sumout ;
wire \hps_0_h2f_axi_master_agent|Add5~9_sumout ;
wire \wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ;
wire \autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ;
wire \link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~4_combout ;
wire \rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ;
wire \data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ;
wire \time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ;
wire \tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ;
wire \spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ;
wire \tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ;
wire \link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ;
wire \hps_0_h2f_axi_master_rd_limiter|has_pending_responses~q ;
wire \router_001|src_data[102]~0_combout ;
wire \hps_0_h2f_axi_master_rd_limiter|last_channel[6]~q ;
wire \router_001|Equal6~0_combout ;
wire \router_001|src_data[100]~1_combout ;
wire \router_001|src_data[101]~2_combout ;
wire \router_001|src_data[103]~3_combout ;
wire \cmd_mux_008|saved_grant[1]~q ;
wire \data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ;
wire \data_o_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \autostart_s1_translator|waitrequest_reset_override~q ;
wire \data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ;
wire \data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ;
wire \data_o_s1_translator|wait_latency_counter[1]~q ;
wire \data_o_s1_translator|wait_latency_counter[0]~q ;
wire \data_o_s1_agent|cp_ready~0_combout ;
wire \data_o_s1_agent|cp_ready~1_combout ;
wire \data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ;
wire \router_001|src_channel~0_combout ;
wire \autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ;
wire \data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ;
wire \data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ;
wire \data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ;
wire \cmd_mux_011|saved_grant[1]~q ;
wire \tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ;
wire \tick_out_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ;
wire \tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ;
wire \tick_out_s1_translator|wait_latency_counter[1]~q ;
wire \tick_out_s1_translator|wait_latency_counter[0]~q ;
wire \tick_out_s1_agent|cp_ready~0_combout ;
wire \tick_out_s1_agent|cp_ready~1_combout ;
wire \tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ;
wire \cmd_mux_011|last_cycle~0_combout ;
wire \tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ;
wire \tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ;
wire \tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ;
wire \cmd_mux_012|saved_grant[1]~q ;
wire \time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ;
wire \time_out_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ;
wire \time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ;
wire \time_out_s1_translator|wait_latency_counter[1]~q ;
wire \time_out_s1_translator|wait_latency_counter[0]~q ;
wire \time_out_s1_agent|cp_ready~0_combout ;
wire \time_out_s1_agent|cp_ready~1_combout ;
wire \time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ;
wire \cmd_mux_012|last_cycle~0_combout ;
wire \time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ;
wire \time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ;
wire \time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ;
wire \link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ;
wire \link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ;
wire \link_disable_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ;
wire \link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ;
wire \link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ;
wire \link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ;
wire \link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ;
wire \link_disable_s1_agent|WideOr0~0_combout ;
wire \link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ;
wire \link_disable_s1_agent|cp_ready~0_combout ;
wire \link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ;
wire \link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ;
wire \cmd_mux_001|saved_grant[1]~q ;
wire \router_001|src_channel[1]~1_combout ;
wire \cmd_demux_001|WideOr0~0_combout ;
wire \tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ;
wire \tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ;
wire \tx_clk_div_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ;
wire \tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ;
wire \tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ;
wire \tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ;
wire \tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ;
wire \tx_clk_div_s1_agent|WideOr0~0_combout ;
wire \tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ;
wire \tx_clk_div_s1_agent|cp_ready~0_combout ;
wire \tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ;
wire \tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ;
wire \cmd_mux_015|saved_grant[1]~q ;
wire \router_001|Equal15~0_combout ;
wire \spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ;
wire \spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ;
wire \spill_enable_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ;
wire \spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ;
wire \spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ;
wire \spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ;
wire \spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ;
wire \spill_enable_s1_agent|WideOr0~0_combout ;
wire \spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ;
wire \spill_enable_s1_agent|cp_ready~0_combout ;
wire \spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ;
wire \spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ;
wire \router_001|Equal16~0_combout ;
wire \cmd_mux_016|saved_grant[1]~q ;
wire \cmd_demux_001|WideOr0~1_combout ;
wire \tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ;
wire \tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ;
wire \tick_in_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ;
wire \tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ;
wire \tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ;
wire \tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ;
wire \tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ;
wire \tick_in_s1_agent|WideOr0~0_combout ;
wire \tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ;
wire \tick_in_s1_agent|cp_ready~0_combout ;
wire \tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ;
wire \tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ;
wire \cmd_mux_013|saved_grant[1]~q ;
wire \router_001|src_channel[13]~2_combout ;
wire \time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ;
wire \time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ;
wire \time_in_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ;
wire \time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ;
wire \time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ;
wire \time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ;
wire \time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ;
wire \time_in_s1_agent|WideOr0~0_combout ;
wire \time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ;
wire \time_in_s1_agent|cp_ready~0_combout ;
wire \time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ;
wire \time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ;
wire \cmd_mux_014|saved_grant[1]~q ;
wire \router_001|Equal14~0_combout ;
wire \cmd_demux_001|WideOr0~2_combout ;
wire \router_001|Equal3~0_combout ;
wire \cmd_mux_003|saved_grant[1]~q ;
wire \currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ;
wire \currentstate_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ;
wire \currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ;
wire \currentstate_s1_translator|wait_latency_counter[1]~q ;
wire \currentstate_s1_translator|wait_latency_counter[0]~q ;
wire \currentstate_s1_agent|cp_ready~0_combout ;
wire \currentstate_s1_agent|cp_ready~1_combout ;
wire \currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ;
wire \currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ;
wire \currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ;
wire \currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ;
wire \data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ;
wire \data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ;
wire \data_i_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ;
wire \data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ;
wire \data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ;
wire \data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ;
wire \data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ;
wire \data_i_s1_agent|WideOr0~0_combout ;
wire \data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ;
wire \data_i_s1_agent|cp_ready~0_combout ;
wire \data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ;
wire \data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ;
wire \cmd_mux_005|saved_grant[1]~q ;
wire \rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ;
wire \rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ;
wire \rd_data_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ;
wire \rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ;
wire \rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ;
wire \rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ;
wire \rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ;
wire \rd_data_s1_agent|WideOr0~0_combout ;
wire \rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ;
wire \rd_data_s1_agent|cp_ready~0_combout ;
wire \rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ;
wire \rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ;
wire \cmd_mux_009|saved_grant[1]~q ;
wire \cmd_mux_010|saved_grant[1]~q ;
wire \router_001|Equal10~0_combout ;
wire \rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ;
wire \rx_empty_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ;
wire \rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ;
wire \rx_empty_s1_translator|wait_latency_counter[1]~q ;
wire \rx_empty_s1_translator|wait_latency_counter[0]~q ;
wire \rx_empty_s1_agent|cp_ready~0_combout ;
wire \rx_empty_s1_agent|cp_ready~1_combout ;
wire \rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ;
wire \rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ;
wire \rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ;
wire \rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ;
wire \cmd_mux|saved_grant[1]~q ;
wire \link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ;
wire \link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ;
wire \link_start_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ;
wire \link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ;
wire \link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ;
wire \link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ;
wire \link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ;
wire \link_start_s1_agent|WideOr0~0_combout ;
wire \link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ;
wire \link_start_s1_agent|cp_ready~0_combout ;
wire \link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ;
wire \link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ;
wire \router_001|src_channel[0]~3_combout ;
wire \flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ;
wire \flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ;
wire \flags_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ;
wire \flags_s1_translator|wait_latency_counter[1]~q ;
wire \flags_s1_translator|wait_latency_counter[0]~q ;
wire \flags_s1_agent|cp_ready~0_combout ;
wire \flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ;
wire \tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ;
wire \tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ;
wire \tx_full_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ;
wire \tx_full_s1_translator|wait_latency_counter[1]~q ;
wire \tx_full_s1_translator|wait_latency_counter[0]~q ;
wire \tx_full_s1_agent|cp_ready~0_combout ;
wire \tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ;
wire \flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ;
wire \flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ;
wire \flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ;
wire \cmd_mux_004|saved_grant[1]~q ;
wire \tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ;
wire \tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ;
wire \tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ;
wire \cmd_mux_007|saved_grant[1]~q ;
wire \autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ;
wire \autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ;
wire \autostart_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ;
wire \autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ;
wire \autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ;
wire \autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ;
wire \autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ;
wire \autostart_s1_agent|WideOr0~0_combout ;
wire \autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ;
wire \autostart_s1_agent|cp_ready~0_combout ;
wire \autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ;
wire \autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ;
wire \cmd_mux_002|saved_grant[1]~q ;
wire \wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ;
wire \wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ;
wire \wr_data_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ;
wire \wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ;
wire \wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ;
wire \wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ;
wire \wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ;
wire \wr_data_s1_agent|WideOr0~0_combout ;
wire \wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ;
wire \wr_data_s1_agent|cp_ready~0_combout ;
wire \wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ;
wire \wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ;
wire \cmd_mux_006|saved_grant[1]~q ;
wire \cmd_demux_001|WideOr0~6_combout ;
wire \hps_0_h2f_axi_master_agent|write_addr_data_both_valid~combout ;
wire \hps_0_h2f_axi_master_wr_limiter|has_pending_responses~q ;
wire \hps_0_h2f_axi_master_agent|sop_enable~q ;
wire \hps_0_h2f_axi_master_agent|align_address_to_size|out_data[8]~0_combout ;
wire \hps_0_h2f_axi_master_agent|align_address_to_size|address_burst[5]~q ;
wire \hps_0_h2f_axi_master_agent|align_address_to_size|out_data[5]~1_combout ;
wire \hps_0_h2f_axi_master_agent|align_address_to_size|address_burst[4]~q ;
wire \hps_0_h2f_axi_master_agent|align_address_to_size|out_data[4]~2_combout ;
wire \hps_0_h2f_axi_master_agent|align_address_to_size|out_data[7]~3_combout ;
wire \hps_0_h2f_axi_master_agent|align_address_to_size|out_data[6]~4_combout ;
wire \router|src_data[102]~0_combout ;
wire \router|Equal5~0_combout ;
wire \router|Equal14~0_combout ;
wire \hps_0_h2f_axi_master_wr_limiter|last_channel[6]~q ;
wire \router|src_data[100]~1_combout ;
wire \router|src_data[101]~2_combout ;
wire \router|Equal16~0_combout ;
wire \router|Equal13~0_combout ;
wire \router|src_data[103]~3_combout ;
wire \router|Equal15~0_combout ;
wire \cmd_mux_015|saved_grant[0]~q ;
wire \router|Equal16~1_combout ;
wire \cmd_mux_016|saved_grant[0]~q ;
wire \cmd_demux|WideOr0~0_combout ;
wire \cmd_mux_013|saved_grant[0]~q ;
wire \cmd_mux_014|saved_grant[0]~q ;
wire \cmd_demux|WideOr0~1_combout ;
wire \cmd_mux_006|saved_grant[0]~q ;
wire \router|Equal9~0_combout ;
wire \cmd_mux_009|saved_grant[0]~q ;
wire \cmd_demux|WideOr0~2_combout ;
wire \cmd_mux|saved_grant[0]~q ;
wire \cmd_mux_001|saved_grant[0]~q ;
wire \cmd_demux|WideOr0~3_combout ;
wire \cmd_mux_002|saved_grant[0]~q ;
wire \cmd_mux_005|saved_grant[0]~q ;
wire \cmd_demux|WideOr0~4_combout ;
wire \cmd_demux|WideOr0~5_combout ;
wire \wr_data_s1_translator|read_latency_shift_reg[0]~q ;
wire \wr_data_s1_agent_rdata_fifo|mem_used[0]~q ;
wire \wr_data_s1_agent_rsp_fifo|mem[0][129]~q ;
wire \wr_data_s1_agent_rsp_fifo|mem_used[0]~q ;
wire \wr_data_s1_agent_rsp_fifo|mem[0][68]~q ;
wire \wr_data_s1_agent_rsp_fifo|mem[0][66]~q ;
wire \rsp_demux_006|src0_valid~combout ;
wire \rd_data_s1_translator|read_latency_shift_reg[0]~q ;
wire \rd_data_s1_agent_rdata_fifo|mem_used[0]~q ;
wire \rd_data_s1_agent_rsp_fifo|mem[0][129]~q ;
wire \rd_data_s1_agent_rsp_fifo|mem_used[0]~q ;
wire \rd_data_s1_agent_rsp_fifo|mem[0][68]~q ;
wire \rd_data_s1_agent_rsp_fifo|mem[0][66]~q ;
wire \rsp_demux_009|src0_valid~combout ;
wire \link_start_s1_translator|read_latency_shift_reg[0]~q ;
wire \link_start_s1_agent_rdata_fifo|mem_used[0]~q ;
wire \link_start_s1_agent_rsp_fifo|mem[0][129]~q ;
wire \link_start_s1_agent_rsp_fifo|mem_used[0]~q ;
wire \link_start_s1_agent_rsp_fifo|mem[0][68]~q ;
wire \link_start_s1_agent_rsp_fifo|mem[0][66]~q ;
wire \rsp_demux|src0_valid~combout ;
wire \link_disable_s1_translator|read_latency_shift_reg[0]~q ;
wire \link_disable_s1_agent_rdata_fifo|mem_used[0]~q ;
wire \link_disable_s1_agent_rsp_fifo|mem[0][129]~q ;
wire \link_disable_s1_agent_rsp_fifo|mem_used[0]~q ;
wire \link_disable_s1_agent_rsp_fifo|mem[0][68]~q ;
wire \link_disable_s1_agent_rsp_fifo|mem[0][66]~q ;
wire \rsp_demux_001|src0_valid~combout ;
wire \autostart_s1_translator|read_latency_shift_reg[0]~q ;
wire \autostart_s1_agent_rdata_fifo|mem_used[0]~q ;
wire \autostart_s1_agent_rsp_fifo|mem[0][129]~q ;
wire \autostart_s1_agent_rsp_fifo|mem_used[0]~q ;
wire \autostart_s1_agent_rsp_fifo|mem[0][68]~q ;
wire \autostart_s1_agent_rsp_fifo|mem[0][66]~q ;
wire \rsp_demux_002|src0_valid~combout ;
wire \data_i_s1_translator|read_latency_shift_reg[0]~q ;
wire \data_i_s1_agent_rdata_fifo|mem_used[0]~q ;
wire \data_i_s1_agent_rsp_fifo|mem[0][129]~q ;
wire \data_i_s1_agent_rsp_fifo|mem_used[0]~q ;
wire \data_i_s1_agent_rsp_fifo|mem[0][68]~q ;
wire \data_i_s1_agent_rsp_fifo|mem[0][66]~q ;
wire \rsp_demux_005|src0_valid~combout ;
wire \tick_in_s1_translator|read_latency_shift_reg[0]~q ;
wire \tick_in_s1_agent_rdata_fifo|mem_used[0]~q ;
wire \tick_in_s1_agent_rsp_fifo|mem[0][129]~q ;
wire \tick_in_s1_agent_rsp_fifo|mem_used[0]~q ;
wire \tick_in_s1_agent_rsp_fifo|mem[0][68]~q ;
wire \tick_in_s1_agent_rsp_fifo|mem[0][66]~q ;
wire \rsp_demux_013|src0_valid~combout ;
wire \time_in_s1_translator|read_latency_shift_reg[0]~q ;
wire \time_in_s1_agent_rdata_fifo|mem_used[0]~q ;
wire \time_in_s1_agent_rsp_fifo|mem[0][129]~q ;
wire \time_in_s1_agent_rsp_fifo|mem_used[0]~q ;
wire \time_in_s1_agent_rsp_fifo|mem[0][68]~q ;
wire \time_in_s1_agent_rsp_fifo|mem[0][66]~q ;
wire \rsp_demux_014|src0_valid~combout ;
wire \tx_clk_div_s1_translator|read_latency_shift_reg[0]~q ;
wire \tx_clk_div_s1_agent_rdata_fifo|mem_used[0]~q ;
wire \tx_clk_div_s1_agent_rsp_fifo|mem[0][129]~q ;
wire \tx_clk_div_s1_agent_rsp_fifo|mem_used[0]~q ;
wire \tx_clk_div_s1_agent_rsp_fifo|mem[0][68]~q ;
wire \tx_clk_div_s1_agent_rsp_fifo|mem[0][66]~q ;
wire \rsp_demux_015|src0_valid~combout ;
wire \spill_enable_s1_translator|read_latency_shift_reg[0]~q ;
wire \spill_enable_s1_agent_rdata_fifo|mem_used[0]~q ;
wire \spill_enable_s1_agent_rsp_fifo|mem[0][129]~q ;
wire \spill_enable_s1_agent_rsp_fifo|mem_used[0]~q ;
wire \spill_enable_s1_agent_rsp_fifo|mem[0][68]~q ;
wire \spill_enable_s1_agent_rsp_fifo|mem[0][66]~q ;
wire \rsp_demux_016|src0_valid~combout ;
wire \spill_enable_s1_agent|comb~0_combout ;
wire \rsp_demux_016|src1_valid~0_combout ;
wire \spill_enable_s1_agent_rsp_fifo|mem[0][130]~q ;
wire \spill_enable_s1_agent|uncompressor|last_packet_beat~0_combout ;
wire \spill_enable_s1_agent_rsp_fifo|mem[0][78]~q ;
wire \spill_enable_s1_agent_rsp_fifo|mem[0][77]~q ;
wire \spill_enable_s1_agent_rsp_fifo|mem[0][76]~q ;
wire \spill_enable_s1_agent_rsp_fifo|mem[0][75]~q ;
wire \spill_enable_s1_agent_rsp_fifo|mem[0][74]~q ;
wire \spill_enable_s1_agent|uncompressor|last_packet_beat~1_combout ;
wire \rsp_mux_001|src_payload~0_combout ;
wire \tx_full_s1_translator|read_latency_shift_reg[0]~q ;
wire \tx_full_s1_agent_rdata_fifo|mem_used[0]~q ;
wire \tx_full_s1_agent_rdata_fifo|empty~combout ;
wire \tx_full_s1_agent_rsp_fifo|mem[0][66]~q ;
wire \tx_full_s1_agent_rsp_fifo|mem_used[0]~q ;
wire \tx_full_s1_agent_rsp_fifo|mem[0][78]~q ;
wire \tx_full_s1_agent_rsp_fifo|mem[0][77]~q ;
wire \tx_full_s1_agent_rsp_fifo|mem[0][76]~q ;
wire \tx_full_s1_agent_rsp_fifo|mem[0][75]~q ;
wire \tx_full_s1_agent_rsp_fifo|mem[0][74]~q ;
wire \tx_full_s1_agent|uncompressor|last_packet_beat~3_combout ;
wire \time_out_s1_agent_rsp_fifo|mem[0][130]~q ;
wire \time_out_s1_translator|read_latency_shift_reg[0]~q ;
wire \time_out_s1_agent_rdata_fifo|mem_used[0]~q ;
wire \time_out_s1_agent_rdata_fifo|empty~combout ;
wire \time_out_s1_agent_rsp_fifo|mem[0][66]~q ;
wire \time_out_s1_agent_rsp_fifo|mem_used[0]~q ;
wire \time_out_s1_agent|uncompressor|last_packet_beat~0_combout ;
wire \time_out_s1_agent_rsp_fifo|mem[0][78]~q ;
wire \time_out_s1_agent_rsp_fifo|mem[0][77]~q ;
wire \time_out_s1_agent_rsp_fifo|mem[0][76]~q ;
wire \time_out_s1_agent_rsp_fifo|mem[0][75]~q ;
wire \time_out_s1_agent_rsp_fifo|mem[0][74]~q ;
wire \time_out_s1_agent|uncompressor|last_packet_beat~1_combout ;
wire \tick_out_s1_agent_rsp_fifo|mem[0][130]~q ;
wire \tick_out_s1_translator|read_latency_shift_reg[0]~q ;
wire \tick_out_s1_agent_rdata_fifo|mem_used[0]~q ;
wire \tick_out_s1_agent_rdata_fifo|empty~combout ;
wire \tick_out_s1_agent_rsp_fifo|mem[0][66]~q ;
wire \tick_out_s1_agent_rsp_fifo|mem_used[0]~q ;
wire \tick_out_s1_agent|uncompressor|last_packet_beat~0_combout ;
wire \tick_out_s1_agent_rsp_fifo|mem[0][78]~q ;
wire \tick_out_s1_agent_rsp_fifo|mem[0][77]~q ;
wire \tick_out_s1_agent_rsp_fifo|mem[0][76]~q ;
wire \tick_out_s1_agent_rsp_fifo|mem[0][75]~q ;
wire \tick_out_s1_agent_rsp_fifo|mem[0][74]~q ;
wire \tick_out_s1_agent|uncompressor|last_packet_beat~1_combout ;
wire \rx_empty_s1_agent_rsp_fifo|mem[0][130]~q ;
wire \rx_empty_s1_translator|read_latency_shift_reg[0]~q ;
wire \rx_empty_s1_agent_rdata_fifo|mem_used[0]~q ;
wire \rx_empty_s1_agent_rdata_fifo|empty~combout ;
wire \rx_empty_s1_agent_rsp_fifo|mem[0][66]~q ;
wire \rx_empty_s1_agent_rsp_fifo|mem_used[0]~q ;
wire \rx_empty_s1_agent|uncompressor|last_packet_beat~0_combout ;
wire \rx_empty_s1_agent_rsp_fifo|mem[0][78]~q ;
wire \rx_empty_s1_agent_rsp_fifo|mem[0][77]~q ;
wire \rx_empty_s1_agent_rsp_fifo|mem[0][76]~q ;
wire \rx_empty_s1_agent_rsp_fifo|mem[0][75]~q ;
wire \rx_empty_s1_agent_rsp_fifo|mem[0][74]~q ;
wire \rx_empty_s1_agent|uncompressor|last_packet_beat~1_combout ;
wire \tx_full_s1_agent_rsp_fifo|mem[0][130]~q ;
wire \data_o_s1_agent_rsp_fifo|mem[0][130]~q ;
wire \data_o_s1_translator|read_latency_shift_reg[0]~q ;
wire \data_o_s1_agent_rdata_fifo|mem_used[0]~q ;
wire \data_o_s1_agent_rdata_fifo|empty~combout ;
wire \data_o_s1_agent_rsp_fifo|mem[0][66]~q ;
wire \data_o_s1_agent_rsp_fifo|mem_used[0]~q ;
wire \data_o_s1_agent|uncompressor|last_packet_beat~0_combout ;
wire \data_o_s1_agent_rsp_fifo|mem[0][78]~q ;
wire \data_o_s1_agent_rsp_fifo|mem[0][77]~q ;
wire \data_o_s1_agent_rsp_fifo|mem[0][76]~q ;
wire \data_o_s1_agent_rsp_fifo|mem[0][75]~q ;
wire \data_o_s1_agent_rsp_fifo|mem[0][74]~q ;
wire \data_o_s1_agent|uncompressor|last_packet_beat~1_combout ;
wire \rsp_mux_001|src_payload[0]~6_combout ;
wire \link_start_s1_agent|comb~0_combout ;
wire \rsp_demux|src1_valid~0_combout ;
wire \link_start_s1_agent_rsp_fifo|mem[0][130]~q ;
wire \link_start_s1_agent|uncompressor|last_packet_beat~0_combout ;
wire \link_start_s1_agent_rsp_fifo|mem[0][78]~q ;
wire \link_start_s1_agent_rsp_fifo|mem[0][77]~q ;
wire \link_start_s1_agent_rsp_fifo|mem[0][76]~q ;
wire \link_start_s1_agent_rsp_fifo|mem[0][75]~q ;
wire \link_start_s1_agent_rsp_fifo|mem[0][74]~q ;
wire \link_start_s1_agent|uncompressor|last_packet_beat~1_combout ;
wire \link_disable_s1_agent|comb~0_combout ;
wire \rsp_demux_001|src1_valid~0_combout ;
wire \link_disable_s1_agent_rsp_fifo|mem[0][130]~q ;
wire \link_disable_s1_agent|uncompressor|last_packet_beat~0_combout ;
wire \link_disable_s1_agent_rsp_fifo|mem[0][78]~q ;
wire \link_disable_s1_agent_rsp_fifo|mem[0][77]~q ;
wire \link_disable_s1_agent_rsp_fifo|mem[0][76]~q ;
wire \link_disable_s1_agent_rsp_fifo|mem[0][75]~q ;
wire \link_disable_s1_agent_rsp_fifo|mem[0][74]~q ;
wire \link_disable_s1_agent|uncompressor|last_packet_beat~1_combout ;
wire \autostart_s1_agent|comb~0_combout ;
wire \rsp_demux_002|src1_valid~0_combout ;
wire \autostart_s1_agent_rsp_fifo|mem[0][130]~q ;
wire \autostart_s1_agent|uncompressor|last_packet_beat~0_combout ;
wire \autostart_s1_agent_rsp_fifo|mem[0][78]~q ;
wire \autostart_s1_agent_rsp_fifo|mem[0][77]~q ;
wire \autostart_s1_agent_rsp_fifo|mem[0][76]~q ;
wire \autostart_s1_agent_rsp_fifo|mem[0][75]~q ;
wire \autostart_s1_agent_rsp_fifo|mem[0][74]~q ;
wire \autostart_s1_agent|uncompressor|last_packet_beat~1_combout ;
wire \data_i_s1_agent|comb~0_combout ;
wire \rsp_demux_005|src1_valid~0_combout ;
wire \data_i_s1_agent_rsp_fifo|mem[0][130]~q ;
wire \data_i_s1_agent|uncompressor|last_packet_beat~0_combout ;
wire \data_i_s1_agent_rsp_fifo|mem[0][78]~q ;
wire \data_i_s1_agent_rsp_fifo|mem[0][77]~q ;
wire \data_i_s1_agent_rsp_fifo|mem[0][76]~q ;
wire \data_i_s1_agent_rsp_fifo|mem[0][75]~q ;
wire \data_i_s1_agent_rsp_fifo|mem[0][74]~q ;
wire \data_i_s1_agent|uncompressor|last_packet_beat~1_combout ;
wire \wr_data_s1_agent|comb~0_combout ;
wire \rsp_demux_006|src1_valid~0_combout ;
wire \wr_data_s1_agent_rsp_fifo|mem[0][130]~q ;
wire \wr_data_s1_agent|uncompressor|last_packet_beat~0_combout ;
wire \wr_data_s1_agent_rsp_fifo|mem[0][78]~q ;
wire \wr_data_s1_agent_rsp_fifo|mem[0][77]~q ;
wire \wr_data_s1_agent_rsp_fifo|mem[0][76]~q ;
wire \wr_data_s1_agent_rsp_fifo|mem[0][75]~q ;
wire \wr_data_s1_agent_rsp_fifo|mem[0][74]~q ;
wire \wr_data_s1_agent|uncompressor|last_packet_beat~1_combout ;
wire \currentstate_s1_agent_rsp_fifo|mem[0][130]~q ;
wire \currentstate_s1_translator|read_latency_shift_reg[0]~q ;
wire \currentstate_s1_agent_rdata_fifo|mem_used[0]~q ;
wire \currentstate_s1_agent_rdata_fifo|empty~combout ;
wire \currentstate_s1_agent_rsp_fifo|mem[0][66]~q ;
wire \currentstate_s1_agent_rsp_fifo|mem_used[0]~q ;
wire \currentstate_s1_agent|uncompressor|last_packet_beat~0_combout ;
wire \currentstate_s1_agent_rsp_fifo|mem[0][78]~q ;
wire \currentstate_s1_agent_rsp_fifo|mem[0][77]~q ;
wire \currentstate_s1_agent_rsp_fifo|mem[0][76]~q ;
wire \currentstate_s1_agent_rsp_fifo|mem[0][75]~q ;
wire \currentstate_s1_agent_rsp_fifo|mem[0][74]~q ;
wire \currentstate_s1_agent|uncompressor|last_packet_beat~1_combout ;
wire \rsp_mux_001|src_payload[0]~13_combout ;
wire \flags_s1_translator|read_latency_shift_reg[0]~q ;
wire \flags_s1_agent_rdata_fifo|mem_used[0]~q ;
wire \flags_s1_agent_rdata_fifo|empty~combout ;
wire \flags_s1_agent_rsp_fifo|mem[0][66]~q ;
wire \flags_s1_agent_rsp_fifo|mem_used[0]~q ;
wire \flags_s1_agent_rsp_fifo|mem[0][78]~q ;
wire \flags_s1_agent_rsp_fifo|mem[0][77]~q ;
wire \flags_s1_agent_rsp_fifo|mem[0][76]~q ;
wire \flags_s1_agent_rsp_fifo|mem[0][75]~q ;
wire \flags_s1_agent_rsp_fifo|mem[0][74]~q ;
wire \flags_s1_agent|uncompressor|last_packet_beat~3_combout ;
wire \rd_data_s1_agent|comb~0_combout ;
wire \rsp_demux_009|src1_valid~0_combout ;
wire \rd_data_s1_agent_rsp_fifo|mem[0][130]~q ;
wire \rd_data_s1_agent|uncompressor|last_packet_beat~0_combout ;
wire \rd_data_s1_agent_rsp_fifo|mem[0][78]~q ;
wire \rd_data_s1_agent_rsp_fifo|mem[0][77]~q ;
wire \rd_data_s1_agent_rsp_fifo|mem[0][76]~q ;
wire \rd_data_s1_agent_rsp_fifo|mem[0][75]~q ;
wire \rd_data_s1_agent_rsp_fifo|mem[0][74]~q ;
wire \rd_data_s1_agent|uncompressor|last_packet_beat~1_combout ;
wire \tick_in_s1_agent|comb~0_combout ;
wire \rsp_demux_013|src1_valid~0_combout ;
wire \tick_in_s1_agent_rsp_fifo|mem[0][130]~q ;
wire \tick_in_s1_agent|uncompressor|last_packet_beat~0_combout ;
wire \tick_in_s1_agent_rsp_fifo|mem[0][78]~q ;
wire \tick_in_s1_agent_rsp_fifo|mem[0][77]~q ;
wire \tick_in_s1_agent_rsp_fifo|mem[0][76]~q ;
wire \tick_in_s1_agent_rsp_fifo|mem[0][75]~q ;
wire \tick_in_s1_agent_rsp_fifo|mem[0][74]~q ;
wire \tick_in_s1_agent|uncompressor|last_packet_beat~1_combout ;
wire \time_in_s1_agent|comb~0_combout ;
wire \rsp_demux_014|src1_valid~0_combout ;
wire \time_in_s1_agent_rsp_fifo|mem[0][130]~q ;
wire \time_in_s1_agent|uncompressor|last_packet_beat~0_combout ;
wire \time_in_s1_agent_rsp_fifo|mem[0][78]~q ;
wire \time_in_s1_agent_rsp_fifo|mem[0][77]~q ;
wire \time_in_s1_agent_rsp_fifo|mem[0][76]~q ;
wire \time_in_s1_agent_rsp_fifo|mem[0][75]~q ;
wire \time_in_s1_agent_rsp_fifo|mem[0][74]~q ;
wire \time_in_s1_agent|uncompressor|last_packet_beat~1_combout ;
wire \tx_clk_div_s1_agent|comb~0_combout ;
wire \rsp_demux_015|src1_valid~0_combout ;
wire \tx_clk_div_s1_agent_rsp_fifo|mem[0][130]~q ;
wire \tx_clk_div_s1_agent|uncompressor|last_packet_beat~0_combout ;
wire \tx_clk_div_s1_agent_rsp_fifo|mem[0][78]~q ;
wire \tx_clk_div_s1_agent_rsp_fifo|mem[0][77]~q ;
wire \tx_clk_div_s1_agent_rsp_fifo|mem[0][76]~q ;
wire \tx_clk_div_s1_agent_rsp_fifo|mem[0][75]~q ;
wire \tx_clk_div_s1_agent_rsp_fifo|mem[0][74]~q ;
wire \tx_clk_div_s1_agent|uncompressor|last_packet_beat~1_combout ;
wire \flags_s1_agent_rsp_fifo|mem[0][130]~q ;
wire \rsp_mux_001|src_payload[0]~19_combout ;
wire \tx_clk_div_s1_agent_rsp_fifo|mem[0][105]~q ;
wire \spill_enable_s1_agent_rsp_fifo|mem[0][105]~q ;
wire \tick_in_s1_agent_rsp_fifo|mem[0][105]~q ;
wire \time_in_s1_agent_rsp_fifo|mem[0][105]~q ;
wire \autostart_s1_agent_rsp_fifo|mem[0][105]~q ;
wire \rd_data_s1_agent_rsp_fifo|mem[0][105]~q ;
wire \link_start_s1_agent_rsp_fifo|mem[0][105]~q ;
wire \link_disable_s1_agent_rsp_fifo|mem[0][105]~q ;
wire \data_i_s1_agent_rsp_fifo|mem[0][105]~q ;
wire \wr_data_s1_agent_rsp_fifo|mem[0][105]~q ;
wire \tx_clk_div_s1_agent_rsp_fifo|mem[0][106]~q ;
wire \spill_enable_s1_agent_rsp_fifo|mem[0][106]~q ;
wire \tick_in_s1_agent_rsp_fifo|mem[0][106]~q ;
wire \time_in_s1_agent_rsp_fifo|mem[0][106]~q ;
wire \autostart_s1_agent_rsp_fifo|mem[0][106]~q ;
wire \rd_data_s1_agent_rsp_fifo|mem[0][106]~q ;
wire \link_start_s1_agent_rsp_fifo|mem[0][106]~q ;
wire \link_disable_s1_agent_rsp_fifo|mem[0][106]~q ;
wire \data_i_s1_agent_rsp_fifo|mem[0][106]~q ;
wire \wr_data_s1_agent_rsp_fifo|mem[0][106]~q ;
wire \tx_clk_div_s1_agent_rsp_fifo|mem[0][107]~q ;
wire \spill_enable_s1_agent_rsp_fifo|mem[0][107]~q ;
wire \tick_in_s1_agent_rsp_fifo|mem[0][107]~q ;
wire \time_in_s1_agent_rsp_fifo|mem[0][107]~q ;
wire \autostart_s1_agent_rsp_fifo|mem[0][107]~q ;
wire \rd_data_s1_agent_rsp_fifo|mem[0][107]~q ;
wire \link_start_s1_agent_rsp_fifo|mem[0][107]~q ;
wire \link_disable_s1_agent_rsp_fifo|mem[0][107]~q ;
wire \data_i_s1_agent_rsp_fifo|mem[0][107]~q ;
wire \wr_data_s1_agent_rsp_fifo|mem[0][107]~q ;
wire \tx_clk_div_s1_agent_rsp_fifo|mem[0][108]~q ;
wire \spill_enable_s1_agent_rsp_fifo|mem[0][108]~q ;
wire \tick_in_s1_agent_rsp_fifo|mem[0][108]~q ;
wire \time_in_s1_agent_rsp_fifo|mem[0][108]~q ;
wire \autostart_s1_agent_rsp_fifo|mem[0][108]~q ;
wire \rd_data_s1_agent_rsp_fifo|mem[0][108]~q ;
wire \link_start_s1_agent_rsp_fifo|mem[0][108]~q ;
wire \link_disable_s1_agent_rsp_fifo|mem[0][108]~q ;
wire \data_i_s1_agent_rsp_fifo|mem[0][108]~q ;
wire \wr_data_s1_agent_rsp_fifo|mem[0][108]~q ;
wire \tx_clk_div_s1_agent_rsp_fifo|mem[0][109]~q ;
wire \spill_enable_s1_agent_rsp_fifo|mem[0][109]~q ;
wire \tick_in_s1_agent_rsp_fifo|mem[0][109]~q ;
wire \time_in_s1_agent_rsp_fifo|mem[0][109]~q ;
wire \autostart_s1_agent_rsp_fifo|mem[0][109]~q ;
wire \rd_data_s1_agent_rsp_fifo|mem[0][109]~q ;
wire \link_start_s1_agent_rsp_fifo|mem[0][109]~q ;
wire \link_disable_s1_agent_rsp_fifo|mem[0][109]~q ;
wire \data_i_s1_agent_rsp_fifo|mem[0][109]~q ;
wire \wr_data_s1_agent_rsp_fifo|mem[0][109]~q ;
wire \tx_clk_div_s1_agent_rsp_fifo|mem[0][110]~q ;
wire \spill_enable_s1_agent_rsp_fifo|mem[0][110]~q ;
wire \tick_in_s1_agent_rsp_fifo|mem[0][110]~q ;
wire \time_in_s1_agent_rsp_fifo|mem[0][110]~q ;
wire \autostart_s1_agent_rsp_fifo|mem[0][110]~q ;
wire \rd_data_s1_agent_rsp_fifo|mem[0][110]~q ;
wire \link_start_s1_agent_rsp_fifo|mem[0][110]~q ;
wire \link_disable_s1_agent_rsp_fifo|mem[0][110]~q ;
wire \data_i_s1_agent_rsp_fifo|mem[0][110]~q ;
wire \wr_data_s1_agent_rsp_fifo|mem[0][110]~q ;
wire \tx_clk_div_s1_agent_rsp_fifo|mem[0][111]~q ;
wire \spill_enable_s1_agent_rsp_fifo|mem[0][111]~q ;
wire \tick_in_s1_agent_rsp_fifo|mem[0][111]~q ;
wire \time_in_s1_agent_rsp_fifo|mem[0][111]~q ;
wire \autostart_s1_agent_rsp_fifo|mem[0][111]~q ;
wire \rd_data_s1_agent_rsp_fifo|mem[0][111]~q ;
wire \link_start_s1_agent_rsp_fifo|mem[0][111]~q ;
wire \link_disable_s1_agent_rsp_fifo|mem[0][111]~q ;
wire \data_i_s1_agent_rsp_fifo|mem[0][111]~q ;
wire \wr_data_s1_agent_rsp_fifo|mem[0][111]~q ;
wire \tx_clk_div_s1_agent_rsp_fifo|mem[0][112]~q ;
wire \spill_enable_s1_agent_rsp_fifo|mem[0][112]~q ;
wire \tick_in_s1_agent_rsp_fifo|mem[0][112]~q ;
wire \time_in_s1_agent_rsp_fifo|mem[0][112]~q ;
wire \autostart_s1_agent_rsp_fifo|mem[0][112]~q ;
wire \rd_data_s1_agent_rsp_fifo|mem[0][112]~q ;
wire \link_start_s1_agent_rsp_fifo|mem[0][112]~q ;
wire \link_disable_s1_agent_rsp_fifo|mem[0][112]~q ;
wire \data_i_s1_agent_rsp_fifo|mem[0][112]~q ;
wire \wr_data_s1_agent_rsp_fifo|mem[0][112]~q ;
wire \tx_clk_div_s1_agent_rsp_fifo|mem[0][113]~q ;
wire \spill_enable_s1_agent_rsp_fifo|mem[0][113]~q ;
wire \tick_in_s1_agent_rsp_fifo|mem[0][113]~q ;
wire \time_in_s1_agent_rsp_fifo|mem[0][113]~q ;
wire \autostart_s1_agent_rsp_fifo|mem[0][113]~q ;
wire \rd_data_s1_agent_rsp_fifo|mem[0][113]~q ;
wire \link_start_s1_agent_rsp_fifo|mem[0][113]~q ;
wire \link_disable_s1_agent_rsp_fifo|mem[0][113]~q ;
wire \data_i_s1_agent_rsp_fifo|mem[0][113]~q ;
wire \wr_data_s1_agent_rsp_fifo|mem[0][113]~q ;
wire \tx_clk_div_s1_agent_rsp_fifo|mem[0][114]~q ;
wire \spill_enable_s1_agent_rsp_fifo|mem[0][114]~q ;
wire \tick_in_s1_agent_rsp_fifo|mem[0][114]~q ;
wire \time_in_s1_agent_rsp_fifo|mem[0][114]~q ;
wire \autostart_s1_agent_rsp_fifo|mem[0][114]~q ;
wire \rd_data_s1_agent_rsp_fifo|mem[0][114]~q ;
wire \link_start_s1_agent_rsp_fifo|mem[0][114]~q ;
wire \link_disable_s1_agent_rsp_fifo|mem[0][114]~q ;
wire \data_i_s1_agent_rsp_fifo|mem[0][114]~q ;
wire \wr_data_s1_agent_rsp_fifo|mem[0][114]~q ;
wire \tx_clk_div_s1_agent_rsp_fifo|mem[0][115]~q ;
wire \spill_enable_s1_agent_rsp_fifo|mem[0][115]~q ;
wire \tick_in_s1_agent_rsp_fifo|mem[0][115]~q ;
wire \time_in_s1_agent_rsp_fifo|mem[0][115]~q ;
wire \autostart_s1_agent_rsp_fifo|mem[0][115]~q ;
wire \rd_data_s1_agent_rsp_fifo|mem[0][115]~q ;
wire \link_start_s1_agent_rsp_fifo|mem[0][115]~q ;
wire \link_disable_s1_agent_rsp_fifo|mem[0][115]~q ;
wire \data_i_s1_agent_rsp_fifo|mem[0][115]~q ;
wire \wr_data_s1_agent_rsp_fifo|mem[0][115]~q ;
wire \tx_clk_div_s1_agent_rsp_fifo|mem[0][116]~q ;
wire \spill_enable_s1_agent_rsp_fifo|mem[0][116]~q ;
wire \tick_in_s1_agent_rsp_fifo|mem[0][116]~q ;
wire \time_in_s1_agent_rsp_fifo|mem[0][116]~q ;
wire \autostart_s1_agent_rsp_fifo|mem[0][116]~q ;
wire \rd_data_s1_agent_rsp_fifo|mem[0][116]~q ;
wire \link_start_s1_agent_rsp_fifo|mem[0][116]~q ;
wire \link_disable_s1_agent_rsp_fifo|mem[0][116]~q ;
wire \data_i_s1_agent_rsp_fifo|mem[0][116]~q ;
wire \wr_data_s1_agent_rsp_fifo|mem[0][116]~q ;
wire \autostart_s1_translator|av_readdata_pre[0]~q ;
wire \autostart_s1_agent_rdata_fifo|mem[0][0]~q ;
wire \tx_clk_div_s1_translator|av_readdata_pre[0]~q ;
wire \tx_clk_div_s1_agent_rdata_fifo|always4~0_combout ;
wire \tx_clk_div_s1_agent_rdata_fifo|mem[0][0]~q ;
wire \currentstate_s1_translator|av_readdata_pre[0]~q ;
wire \data_o_s1_translator|av_readdata_pre[0]~q ;
wire \tx_full_s1_agent_rdata_fifo|mem[0][0]~q ;
wire \tx_full_s1_translator|av_readdata_pre[0]~q ;
wire \flags_s1_translator|av_readdata_pre[0]~q ;
wire \flags_s1_agent_rdata_fifo|mem[0][0]~q ;
wire \time_out_s1_agent_rdata_fifo|mem[0][0]~q ;
wire \time_out_s1_translator|av_readdata_pre[0]~q ;
wire \data_o_s1_agent_rdata_fifo|mem[0][0]~q ;
wire \tick_out_s1_translator|av_readdata_pre[0]~q ;
wire \tick_out_s1_agent_rdata_fifo|mem[0][0]~q ;
wire \rx_empty_s1_translator|av_readdata_pre[0]~q ;
wire \currentstate_s1_agent_rdata_fifo|mem[0][0]~q ;
wire \rx_empty_s1_agent_rdata_fifo|mem[0][0]~q ;
wire \link_start_s1_translator|av_readdata_pre[0]~q ;
wire \link_start_s1_agent_rdata_fifo|mem[0][0]~q ;
wire \link_disable_s1_translator|av_readdata_pre[0]~q ;
wire \link_disable_s1_agent_rdata_fifo|mem[0][0]~q ;
wire \wr_data_s1_translator|av_readdata_pre[0]~q ;
wire \wr_data_s1_agent_rdata_fifo|mem[0][0]~q ;
wire \rd_data_s1_translator|av_readdata_pre[0]~q ;
wire \rd_data_s1_agent_rdata_fifo|mem[0][0]~q ;
wire \tick_in_s1_translator|av_readdata_pre[0]~q ;
wire \tick_in_s1_agent_rdata_fifo|mem[0][0]~q ;
wire \spill_enable_s1_translator|av_readdata_pre[0]~q ;
wire \spill_enable_s1_agent_rdata_fifo|mem[0][0]~q ;
wire \data_i_s1_translator|av_readdata_pre[0]~q ;
wire \data_i_s1_agent_rdata_fifo|always4~0_combout ;
wire \data_i_s1_agent_rdata_fifo|mem[0][0]~q ;
wire \time_in_s1_translator|av_readdata_pre[0]~q ;
wire \time_in_s1_agent_rdata_fifo|always4~0_combout ;
wire \time_in_s1_agent_rdata_fifo|mem[0][0]~q ;
wire \currentstate_s1_translator|av_readdata_pre[1]~q ;
wire \data_i_s1_translator|av_readdata_pre[1]~q ;
wire \data_i_s1_agent_rdata_fifo|mem[0][1]~q ;
wire \data_o_s1_agent_rdata_fifo|mem[0][1]~q ;
wire \time_out_s1_agent_rdata_fifo|mem[0][1]~q ;
wire \time_out_s1_translator|av_readdata_pre[1]~q ;
wire \data_o_s1_translator|av_readdata_pre[1]~q ;
wire \flags_s1_agent_rdata_fifo|mem[0][1]~q ;
wire \flags_s1_translator|av_readdata_pre[1]~q ;
wire \currentstate_s1_agent_rdata_fifo|mem[0][1]~q ;
wire \time_in_s1_translator|av_readdata_pre[1]~q ;
wire \time_in_s1_agent_rdata_fifo|mem[0][1]~q ;
wire \tx_clk_div_s1_translator|av_readdata_pre[1]~q ;
wire \tx_clk_div_s1_agent_rdata_fifo|mem[0][1]~q ;
wire \currentstate_s1_translator|av_readdata_pre[2]~q ;
wire \data_i_s1_translator|av_readdata_pre[2]~q ;
wire \data_i_s1_agent_rdata_fifo|mem[0][2]~q ;
wire \data_o_s1_agent_rdata_fifo|mem[0][2]~q ;
wire \time_out_s1_agent_rdata_fifo|mem[0][2]~q ;
wire \time_out_s1_translator|av_readdata_pre[2]~q ;
wire \data_o_s1_translator|av_readdata_pre[2]~q ;
wire \flags_s1_agent_rdata_fifo|mem[0][2]~q ;
wire \flags_s1_translator|av_readdata_pre[2]~q ;
wire \currentstate_s1_agent_rdata_fifo|mem[0][2]~q ;
wire \time_in_s1_translator|av_readdata_pre[2]~q ;
wire \time_in_s1_agent_rdata_fifo|mem[0][2]~q ;
wire \tx_clk_div_s1_translator|av_readdata_pre[2]~q ;
wire \tx_clk_div_s1_agent_rdata_fifo|mem[0][2]~q ;
wire \flags_s1_translator|av_readdata_pre[3]~q ;
wire \data_i_s1_translator|av_readdata_pre[3]~q ;
wire \data_i_s1_agent_rdata_fifo|mem[0][3]~q ;
wire \data_o_s1_agent_rdata_fifo|mem[0][3]~q ;
wire \time_out_s1_agent_rdata_fifo|mem[0][3]~q ;
wire \time_out_s1_translator|av_readdata_pre[3]~q ;
wire \data_o_s1_translator|av_readdata_pre[3]~q ;
wire \flags_s1_agent_rdata_fifo|mem[0][3]~q ;
wire \time_in_s1_translator|av_readdata_pre[3]~q ;
wire \time_in_s1_agent_rdata_fifo|mem[0][3]~q ;
wire \tx_clk_div_s1_translator|av_readdata_pre[3]~q ;
wire \tx_clk_div_s1_agent_rdata_fifo|mem[0][3]~q ;
wire \flags_s1_translator|av_readdata_pre[4]~q ;
wire \data_i_s1_translator|av_readdata_pre[4]~q ;
wire \data_i_s1_agent_rdata_fifo|mem[0][4]~q ;
wire \data_o_s1_agent_rdata_fifo|mem[0][4]~q ;
wire \time_out_s1_agent_rdata_fifo|mem[0][4]~q ;
wire \time_out_s1_translator|av_readdata_pre[4]~q ;
wire \data_o_s1_translator|av_readdata_pre[4]~q ;
wire \flags_s1_agent_rdata_fifo|mem[0][4]~q ;
wire \time_in_s1_translator|av_readdata_pre[4]~q ;
wire \time_in_s1_agent_rdata_fifo|mem[0][4]~q ;
wire \tx_clk_div_s1_translator|av_readdata_pre[4]~q ;
wire \tx_clk_div_s1_agent_rdata_fifo|mem[0][4]~q ;
wire \flags_s1_translator|av_readdata_pre[5]~q ;
wire \data_i_s1_translator|av_readdata_pre[5]~q ;
wire \data_i_s1_agent_rdata_fifo|mem[0][5]~q ;
wire \data_o_s1_agent_rdata_fifo|mem[0][5]~q ;
wire \time_out_s1_agent_rdata_fifo|mem[0][5]~q ;
wire \time_out_s1_translator|av_readdata_pre[5]~q ;
wire \data_o_s1_translator|av_readdata_pre[5]~q ;
wire \flags_s1_agent_rdata_fifo|mem[0][5]~q ;
wire \time_in_s1_translator|av_readdata_pre[5]~q ;
wire \time_in_s1_agent_rdata_fifo|mem[0][5]~q ;
wire \tx_clk_div_s1_translator|av_readdata_pre[5]~q ;
wire \tx_clk_div_s1_agent_rdata_fifo|mem[0][5]~q ;
wire \flags_s1_translator|av_readdata_pre[6]~q ;
wire \data_i_s1_translator|av_readdata_pre[6]~q ;
wire \data_i_s1_agent_rdata_fifo|mem[0][6]~q ;
wire \data_o_s1_agent_rdata_fifo|mem[0][6]~q ;
wire \time_out_s1_agent_rdata_fifo|mem[0][6]~q ;
wire \time_out_s1_translator|av_readdata_pre[6]~q ;
wire \data_o_s1_translator|av_readdata_pre[6]~q ;
wire \flags_s1_agent_rdata_fifo|mem[0][6]~q ;
wire \time_in_s1_translator|av_readdata_pre[6]~q ;
wire \time_in_s1_agent_rdata_fifo|mem[0][6]~q ;
wire \tx_clk_div_s1_translator|av_readdata_pre[6]~q ;
wire \tx_clk_div_s1_agent_rdata_fifo|mem[0][6]~q ;
wire \flags_s1_translator|av_readdata_pre[7]~q ;
wire \data_i_s1_translator|av_readdata_pre[7]~q ;
wire \data_i_s1_agent_rdata_fifo|mem[0][7]~q ;
wire \time_in_s1_translator|av_readdata_pre[7]~q ;
wire \time_in_s1_agent_rdata_fifo|mem[0][7]~q ;
wire \data_o_s1_agent_rdata_fifo|mem[0][7]~q ;
wire \time_out_s1_agent_rdata_fifo|mem[0][7]~q ;
wire \time_out_s1_translator|av_readdata_pre[7]~q ;
wire \data_o_s1_translator|av_readdata_pre[7]~q ;
wire \flags_s1_agent_rdata_fifo|mem[0][7]~q ;
wire \data_i_s1_translator|av_readdata_pre[8]~q ;
wire \data_i_s1_agent_rdata_fifo|mem[0][8]~q ;
wire \flags_s1_agent_rdata_fifo|mem[0][8]~q ;
wire \flags_s1_translator|av_readdata_pre[8]~q ;
wire \data_o_s1_agent_rdata_fifo|mem[0][8]~q ;
wire \data_o_s1_translator|av_readdata_pre[8]~q ;
wire \flags_s1_agent_rdata_fifo|mem[0][9]~q ;
wire \flags_s1_translator|av_readdata_pre[9]~q ;
wire \flags_s1_agent_rdata_fifo|mem[0][10]~q ;
wire \flags_s1_translator|av_readdata_pre[10]~q ;
wire \time_out_s1_agent_rsp_fifo|mem[0][105]~q ;
wire \currentstate_s1_agent_rsp_fifo|mem[0][105]~q ;
wire \flags_s1_agent_rsp_fifo|mem[0][105]~q ;
wire \tx_full_s1_agent_rsp_fifo|mem[0][105]~q ;
wire \data_o_s1_agent_rsp_fifo|mem[0][105]~q ;
wire \rx_empty_s1_agent_rsp_fifo|mem[0][105]~q ;
wire \tick_out_s1_agent_rsp_fifo|mem[0][105]~q ;
wire \time_out_s1_agent_rsp_fifo|mem[0][106]~q ;
wire \currentstate_s1_agent_rsp_fifo|mem[0][106]~q ;
wire \flags_s1_agent_rsp_fifo|mem[0][106]~q ;
wire \tx_full_s1_agent_rsp_fifo|mem[0][106]~q ;
wire \data_o_s1_agent_rsp_fifo|mem[0][106]~q ;
wire \rx_empty_s1_agent_rsp_fifo|mem[0][106]~q ;
wire \tick_out_s1_agent_rsp_fifo|mem[0][106]~q ;
wire \time_out_s1_agent_rsp_fifo|mem[0][107]~q ;
wire \currentstate_s1_agent_rsp_fifo|mem[0][107]~q ;
wire \flags_s1_agent_rsp_fifo|mem[0][107]~q ;
wire \tx_full_s1_agent_rsp_fifo|mem[0][107]~q ;
wire \data_o_s1_agent_rsp_fifo|mem[0][107]~q ;
wire \rx_empty_s1_agent_rsp_fifo|mem[0][107]~q ;
wire \tick_out_s1_agent_rsp_fifo|mem[0][107]~q ;
wire \time_out_s1_agent_rsp_fifo|mem[0][108]~q ;
wire \currentstate_s1_agent_rsp_fifo|mem[0][108]~q ;
wire \flags_s1_agent_rsp_fifo|mem[0][108]~q ;
wire \tx_full_s1_agent_rsp_fifo|mem[0][108]~q ;
wire \data_o_s1_agent_rsp_fifo|mem[0][108]~q ;
wire \rx_empty_s1_agent_rsp_fifo|mem[0][108]~q ;
wire \tick_out_s1_agent_rsp_fifo|mem[0][108]~q ;
wire \time_out_s1_agent_rsp_fifo|mem[0][109]~q ;
wire \currentstate_s1_agent_rsp_fifo|mem[0][109]~q ;
wire \flags_s1_agent_rsp_fifo|mem[0][109]~q ;
wire \tx_full_s1_agent_rsp_fifo|mem[0][109]~q ;
wire \data_o_s1_agent_rsp_fifo|mem[0][109]~q ;
wire \rx_empty_s1_agent_rsp_fifo|mem[0][109]~q ;
wire \tick_out_s1_agent_rsp_fifo|mem[0][109]~q ;
wire \time_out_s1_agent_rsp_fifo|mem[0][110]~q ;
wire \currentstate_s1_agent_rsp_fifo|mem[0][110]~q ;
wire \flags_s1_agent_rsp_fifo|mem[0][110]~q ;
wire \tx_full_s1_agent_rsp_fifo|mem[0][110]~q ;
wire \data_o_s1_agent_rsp_fifo|mem[0][110]~q ;
wire \rx_empty_s1_agent_rsp_fifo|mem[0][110]~q ;
wire \tick_out_s1_agent_rsp_fifo|mem[0][110]~q ;
wire \time_out_s1_agent_rsp_fifo|mem[0][111]~q ;
wire \currentstate_s1_agent_rsp_fifo|mem[0][111]~q ;
wire \flags_s1_agent_rsp_fifo|mem[0][111]~q ;
wire \tx_full_s1_agent_rsp_fifo|mem[0][111]~q ;
wire \data_o_s1_agent_rsp_fifo|mem[0][111]~q ;
wire \rx_empty_s1_agent_rsp_fifo|mem[0][111]~q ;
wire \tick_out_s1_agent_rsp_fifo|mem[0][111]~q ;
wire \time_out_s1_agent_rsp_fifo|mem[0][112]~q ;
wire \currentstate_s1_agent_rsp_fifo|mem[0][112]~q ;
wire \flags_s1_agent_rsp_fifo|mem[0][112]~q ;
wire \tx_full_s1_agent_rsp_fifo|mem[0][112]~q ;
wire \data_o_s1_agent_rsp_fifo|mem[0][112]~q ;
wire \rx_empty_s1_agent_rsp_fifo|mem[0][112]~q ;
wire \tick_out_s1_agent_rsp_fifo|mem[0][112]~q ;
wire \time_out_s1_agent_rsp_fifo|mem[0][113]~q ;
wire \currentstate_s1_agent_rsp_fifo|mem[0][113]~q ;
wire \flags_s1_agent_rsp_fifo|mem[0][113]~q ;
wire \tx_full_s1_agent_rsp_fifo|mem[0][113]~q ;
wire \data_o_s1_agent_rsp_fifo|mem[0][113]~q ;
wire \rx_empty_s1_agent_rsp_fifo|mem[0][113]~q ;
wire \tick_out_s1_agent_rsp_fifo|mem[0][113]~q ;
wire \time_out_s1_agent_rsp_fifo|mem[0][114]~q ;
wire \currentstate_s1_agent_rsp_fifo|mem[0][114]~q ;
wire \flags_s1_agent_rsp_fifo|mem[0][114]~q ;
wire \tx_full_s1_agent_rsp_fifo|mem[0][114]~q ;
wire \data_o_s1_agent_rsp_fifo|mem[0][114]~q ;
wire \rx_empty_s1_agent_rsp_fifo|mem[0][114]~q ;
wire \tick_out_s1_agent_rsp_fifo|mem[0][114]~q ;
wire \time_out_s1_agent_rsp_fifo|mem[0][115]~q ;
wire \currentstate_s1_agent_rsp_fifo|mem[0][115]~q ;
wire \flags_s1_agent_rsp_fifo|mem[0][115]~q ;
wire \tx_full_s1_agent_rsp_fifo|mem[0][115]~q ;
wire \data_o_s1_agent_rsp_fifo|mem[0][115]~q ;
wire \rx_empty_s1_agent_rsp_fifo|mem[0][115]~q ;
wire \tick_out_s1_agent_rsp_fifo|mem[0][115]~q ;
wire \time_out_s1_agent_rsp_fifo|mem[0][116]~q ;
wire \currentstate_s1_agent_rsp_fifo|mem[0][116]~q ;
wire \flags_s1_agent_rsp_fifo|mem[0][116]~q ;
wire \tx_full_s1_agent_rsp_fifo|mem[0][116]~q ;
wire \data_o_s1_agent_rsp_fifo|mem[0][116]~q ;
wire \rx_empty_s1_agent_rsp_fifo|mem[0][116]~q ;
wire \tick_out_s1_agent_rsp_fifo|mem[0][116]~q ;
wire \data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ;
wire \hps_0_h2f_axi_master_rd_limiter|last_channel[8]~q ;
wire \cmd_mux_008|src_valid~0_combout ;
wire \data_o_s1_agent|uncompressor|last_packet_beat~2_combout ;
wire \data_o_s1_agent_rsp_fifo|write~0_combout ;
wire \data_o_s1_agent_rsp_fifo|write~1_combout ;
wire \hps_0_h2f_axi_master_agent|Decoder1~0_combout ;
wire \data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ;
wire \hps_0_h2f_axi_master_agent|Add2~0_combout ;
wire \hps_0_h2f_axi_master_agent|Add2~1_combout ;
wire \hps_0_h2f_axi_master_agent|Add2~2_combout ;
wire \hps_0_h2f_axi_master_agent|Add2~3_combout ;
wire \data_o_s1_agent|cp_ready~2_combout ;
wire \data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ;
wire \data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ;
wire \data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ;
wire \data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ;
wire \data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ;
wire \tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ;
wire \hps_0_h2f_axi_master_rd_limiter|last_channel[11]~q ;
wire \cmd_mux_011|src_valid~0_combout ;
wire \tick_out_s1_agent|uncompressor|last_packet_beat~2_combout ;
wire \tick_out_s1_agent_rsp_fifo|write~0_combout ;
wire \tick_out_s1_agent_rsp_fifo|write~1_combout ;
wire \tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ;
wire \tick_out_s1_agent|cp_ready~2_combout ;
wire \tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ;
wire \tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ;
wire \tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ;
wire \tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ;
wire \tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ;
wire \time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ;
wire \hps_0_h2f_axi_master_rd_limiter|last_channel[12]~q ;
wire \cmd_mux_012|src_valid~0_combout ;
wire \time_out_s1_agent|uncompressor|last_packet_beat~2_combout ;
wire \time_out_s1_agent_rsp_fifo|write~0_combout ;
wire \time_out_s1_agent_rsp_fifo|write~1_combout ;
wire \time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ;
wire \time_out_s1_agent|cp_ready~2_combout ;
wire \time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ;
wire \time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ;
wire \time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ;
wire \time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ;
wire \time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ;
wire \link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ;
wire \router|Equal5~1_combout ;
wire \hps_0_h2f_axi_master_wr_limiter|last_channel[1]~q ;
wire \cmd_demux|src1_valid~0_combout ;
wire \cmd_demux|src1_valid~1_combout ;
wire \hps_0_h2f_axi_master_rd_limiter|last_channel[1]~q ;
wire \cmd_mux_001|src_valid~0_combout ;
wire \link_disable_s1_agent|cp_ready~3_combout ;
wire \link_disable_s1_agent|uncompressor|last_packet_beat~2_combout ;
wire \rsp_demux_001|WideOr0~0_combout ;
wire \link_disable_s1_agent_rsp_fifo|read~0_combout ;
wire \link_disable_s1_agent|cp_ready~4_combout ;
wire \link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ;
wire \link_disable_s1_agent|rf_source_valid~0_combout ;
wire \cmd_mux_001|src_data[87]~combout ;
wire \cmd_mux_001|src_data[88]~combout ;
wire \cmd_mux_001|src_valid~1_combout ;
wire \cmd_mux_001|src_data[35]~combout ;
wire \cmd_mux_001|src_data[34]~combout ;
wire \cmd_mux_001|src_data[33]~combout ;
wire \cmd_mux_001|src_data[32]~combout ;
wire \link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ;
wire \link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ;
wire \link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ;
wire \link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ;
wire \link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ;
wire \link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ;
wire \cmd_mux_001|src_payload[0]~combout ;
wire \cmd_demux|src1_valid~2_combout ;
wire \hps_0_h2f_axi_master_agent|burst_bytecount[5]~q ;
wire \hps_0_h2f_axi_master_agent|write_cp_data[77]~0_combout ;
wire \hps_0_h2f_axi_master_agent|burst_bytecount[6]~q ;
wire \hps_0_h2f_axi_master_agent|write_cp_data[78]~1_combout ;
wire \hps_0_h2f_axi_master_agent|burst_bytecount[3]~q ;
wire \hps_0_h2f_axi_master_agent|write_cp_data[75]~2_combout ;
wire \hps_0_h2f_axi_master_agent|burst_bytecount[2]~q ;
wire \hps_0_h2f_axi_master_agent|write_cp_data[74]~3_combout ;
wire \hps_0_h2f_axi_master_agent|burst_bytecount[4]~q ;
wire \hps_0_h2f_axi_master_agent|write_cp_data[76]~4_combout ;
wire \link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|WideNor0~0_combout ;
wire \cmd_demux_001|src1_valid~0_combout ;
wire \tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ;
wire \router|Equal15~1_combout ;
wire \hps_0_h2f_axi_master_wr_limiter|last_channel[15]~q ;
wire \cmd_demux|src15_valid~0_combout ;
wire \cmd_demux|src15_valid~1_combout ;
wire \hps_0_h2f_axi_master_rd_limiter|last_channel[15]~q ;
wire \cmd_demux_001|src15_valid~0_combout ;
wire \cmd_mux_015|src_valid~0_combout ;
wire \tx_clk_div_s1_agent|cp_ready~3_combout ;
wire \tx_clk_div_s1_agent|uncompressor|last_packet_beat~2_combout ;
wire \rsp_demux_015|WideOr0~0_combout ;
wire \tx_clk_div_s1_agent_rsp_fifo|read~0_combout ;
wire \tx_clk_div_s1_agent|cp_ready~4_combout ;
wire \tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ;
wire \tx_clk_div_s1_agent|rf_source_valid~0_combout ;
wire \cmd_mux_015|src_data[87]~combout ;
wire \cmd_mux_015|src_data[88]~combout ;
wire \cmd_mux_015|src_valid~1_combout ;
wire \cmd_mux_015|src_data[35]~combout ;
wire \cmd_mux_015|src_data[34]~combout ;
wire \cmd_mux_015|src_data[33]~combout ;
wire \cmd_mux_015|src_data[32]~combout ;
wire \tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ;
wire \tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ;
wire \tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ;
wire \tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ;
wire \tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ;
wire \tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ;
wire \cmd_mux_015|src_payload[0]~combout ;
wire \cmd_demux|src15_valid~2_combout ;
wire \cmd_demux_001|src15_valid~1_combout ;
wire \spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ;
wire \hps_0_h2f_axi_master_wr_limiter|last_channel[16]~q ;
wire \cmd_demux|src16_valid~0_combout ;
wire \cmd_demux|src16_valid~1_combout ;
wire \hps_0_h2f_axi_master_rd_limiter|last_channel[16]~q ;
wire \cmd_demux_001|src16_valid~0_combout ;
wire \cmd_mux_016|src_valid~0_combout ;
wire \cmd_mux_016|src_valid~1_combout ;
wire \cmd_demux|src16_valid~2_combout ;
wire \cmd_mux_016|WideOr1~combout ;
wire \spill_enable_s1_agent|cp_ready~1_combout ;
wire \spill_enable_s1_agent|cp_ready~2_combout ;
wire \spill_enable_s1_agent|uncompressor|last_packet_beat~2_combout ;
wire \rsp_demux_016|WideOr0~0_combout ;
wire \spill_enable_s1_agent_rsp_fifo|read~0_combout ;
wire \spill_enable_s1_agent|cp_ready~3_combout ;
wire \spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ;
wire \spill_enable_s1_agent|rf_source_valid~0_combout ;
wire \cmd_mux_016|src_data[87]~combout ;
wire \cmd_mux_016|src_data[88]~combout ;
wire \cmd_mux_016|src_data[35]~combout ;
wire \cmd_mux_016|src_data[34]~combout ;
wire \cmd_mux_016|src_data[33]~combout ;
wire \cmd_mux_016|src_data[32]~combout ;
wire \spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ;
wire \spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ;
wire \spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ;
wire \spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ;
wire \spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ;
wire \spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ;
wire \cmd_mux_016|src_payload[0]~combout ;
wire \cmd_demux_001|src16_valid~1_combout ;
wire \tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ;
wire \hps_0_h2f_axi_master_wr_limiter|last_channel[13]~q ;
wire \cmd_demux|src13_valid~0_combout ;
wire \cmd_demux|src13_valid~1_combout ;
wire \hps_0_h2f_axi_master_rd_limiter|last_channel[13]~q ;
wire \cmd_mux_013|src_valid~2_combout ;
wire \tick_in_s1_agent|cp_ready~3_combout ;
wire \tick_in_s1_agent|uncompressor|last_packet_beat~2_combout ;
wire \rsp_demux_013|WideOr0~0_combout ;
wire \tick_in_s1_agent_rsp_fifo|read~0_combout ;
wire \tick_in_s1_agent|cp_ready~4_combout ;
wire \tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ;
wire \tick_in_s1_agent|rf_source_valid~0_combout ;
wire \cmd_mux_013|src_data[87]~combout ;
wire \cmd_mux_013|src_data[88]~combout ;
wire \cmd_mux_013|src_valid~3_combout ;
wire \cmd_mux_013|src_data[35]~combout ;
wire \cmd_mux_013|src_data[34]~combout ;
wire \cmd_mux_013|src_data[33]~combout ;
wire \cmd_mux_013|src_data[32]~combout ;
wire \tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ;
wire \tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ;
wire \tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ;
wire \tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ;
wire \tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ;
wire \tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ;
wire \cmd_mux_013|src_payload[0]~combout ;
wire \cmd_demux|src13_valid~2_combout ;
wire \time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ;
wire \router|Equal14~1_combout ;
wire \hps_0_h2f_axi_master_wr_limiter|last_channel[14]~q ;
wire \cmd_demux|src14_valid~0_combout ;
wire \cmd_demux|src14_valid~1_combout ;
wire \hps_0_h2f_axi_master_rd_limiter|last_channel[14]~q ;
wire \cmd_demux_001|src14_valid~0_combout ;
wire \cmd_mux_014|src_valid~0_combout ;
wire \time_in_s1_agent|cp_ready~3_combout ;
wire \time_in_s1_agent|uncompressor|last_packet_beat~2_combout ;
wire \rsp_demux_014|WideOr0~0_combout ;
wire \time_in_s1_agent_rsp_fifo|read~0_combout ;
wire \time_in_s1_agent|cp_ready~4_combout ;
wire \time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ;
wire \time_in_s1_agent|rf_source_valid~0_combout ;
wire \cmd_mux_014|src_data[87]~combout ;
wire \cmd_mux_014|src_data[88]~combout ;
wire \cmd_mux_014|src_valid~1_combout ;
wire \cmd_mux_014|src_data[35]~combout ;
wire \cmd_mux_014|src_data[34]~combout ;
wire \cmd_mux_014|src_data[33]~combout ;
wire \cmd_mux_014|src_data[32]~combout ;
wire \time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ;
wire \time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ;
wire \time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ;
wire \time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ;
wire \time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ;
wire \time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ;
wire \cmd_mux_014|src_payload[0]~combout ;
wire \cmd_demux|src14_valid~2_combout ;
wire \cmd_demux_001|src14_valid~1_combout ;
wire \currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ;
wire \hps_0_h2f_axi_master_rd_limiter|last_channel[3]~q ;
wire \cmd_mux_003|src_valid~0_combout ;
wire \currentstate_s1_agent|uncompressor|last_packet_beat~2_combout ;
wire \currentstate_s1_agent_rsp_fifo|write~0_combout ;
wire \currentstate_s1_agent_rsp_fifo|write~1_combout ;
wire \currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ;
wire \currentstate_s1_agent|cp_ready~2_combout ;
wire \currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ;
wire \currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ;
wire \currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ;
wire \currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ;
wire \currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ;
wire \data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ;
wire \hps_0_h2f_axi_master_wr_limiter|last_channel[5]~q ;
wire \cmd_demux|src5_valid~0_combout ;
wire \cmd_demux|src5_valid~1_combout ;
wire \hps_0_h2f_axi_master_rd_limiter|cmd_src_valid[5]~0_combout ;
wire \cmd_mux_005|src_valid~1_combout ;
wire \data_i_s1_agent|cp_ready~3_combout ;
wire \data_i_s1_agent|uncompressor|last_packet_beat~2_combout ;
wire \rsp_demux_005|WideOr0~0_combout ;
wire \data_i_s1_agent_rsp_fifo|read~0_combout ;
wire \data_i_s1_agent|cp_ready~4_combout ;
wire \data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ;
wire \data_i_s1_agent|rf_source_valid~0_combout ;
wire \cmd_mux_005|src_data[87]~combout ;
wire \cmd_mux_005|src_data[88]~combout ;
wire \cmd_mux_005|src_valid~2_combout ;
wire \cmd_mux_005|src_data[35]~combout ;
wire \cmd_mux_005|src_data[34]~combout ;
wire \cmd_mux_005|src_data[33]~combout ;
wire \cmd_mux_005|src_data[32]~combout ;
wire \data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ;
wire \data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ;
wire \data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ;
wire \data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ;
wire \data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ;
wire \data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ;
wire \cmd_mux_005|src_payload[0]~combout ;
wire \cmd_demux|src5_valid~2_combout ;
wire \rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ;
wire \hps_0_h2f_axi_master_wr_limiter|last_channel[9]~q ;
wire \cmd_demux|src9_valid~0_combout ;
wire \cmd_demux|src9_valid~1_combout ;
wire \router_001|Equal9~0_combout ;
wire \hps_0_h2f_axi_master_rd_limiter|last_channel[9]~q ;
wire \cmd_demux_001|src9_valid~0_combout ;
wire \cmd_mux_009|src_valid~0_combout ;
wire \rd_data_s1_agent|cp_ready~3_combout ;
wire \rd_data_s1_agent|uncompressor|last_packet_beat~2_combout ;
wire \rsp_demux_009|WideOr0~0_combout ;
wire \rd_data_s1_agent_rsp_fifo|read~0_combout ;
wire \rd_data_s1_agent|cp_ready~4_combout ;
wire \rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ;
wire \rd_data_s1_agent|rf_source_valid~0_combout ;
wire \cmd_mux_009|src_data[87]~combout ;
wire \cmd_mux_009|src_data[88]~combout ;
wire \cmd_mux_009|src_valid~1_combout ;
wire \cmd_mux_009|src_data[35]~combout ;
wire \cmd_mux_009|src_data[34]~combout ;
wire \cmd_mux_009|src_data[33]~combout ;
wire \cmd_mux_009|src_data[32]~combout ;
wire \rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ;
wire \rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ;
wire \rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ;
wire \rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ;
wire \rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ;
wire \rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ;
wire \cmd_mux_009|src_payload[0]~combout ;
wire \cmd_demux|src9_valid~2_combout ;
wire \cmd_demux_001|src9_valid~1_combout ;
wire \hps_0_h2f_axi_master_rd_limiter|last_channel[10]~q ;
wire \cmd_mux_010|src_valid~0_combout ;
wire \rx_empty_s1_agent|uncompressor|last_packet_beat~2_combout ;
wire \rx_empty_s1_agent_rsp_fifo|write~0_combout ;
wire \rx_empty_s1_agent_rsp_fifo|write~1_combout ;
wire \rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ;
wire \rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ;
wire \rx_empty_s1_agent|cp_ready~2_combout ;
wire \rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ;
wire \rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ;
wire \rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ;
wire \rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ;
wire \rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ;
wire \hps_0_h2f_axi_master_wr_limiter|last_channel[0]~q ;
wire \cmd_demux|src0_valid~1_combout ;
wire \hps_0_h2f_axi_master_rd_limiter|last_channel[0]~q ;
wire \cmd_demux_001|src0_valid~0_combout ;
wire \link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ;
wire \cmd_mux|src_valid~0_combout ;
wire \cmd_mux|src_payload[0]~combout ;
wire \link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ;
wire \link_start_s1_agent|cp_ready~2_combout ;
wire \link_start_s1_agent|uncompressor|last_packet_beat~2_combout ;
wire \rsp_demux|WideOr0~0_combout ;
wire \link_start_s1_agent_rsp_fifo|read~0_combout ;
wire \link_start_s1_agent|cp_ready~3_combout ;
wire \link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ;
wire \link_start_s1_agent|rf_source_valid~0_combout ;
wire \cmd_mux|src_data[87]~combout ;
wire \cmd_mux|src_data[88]~combout ;
wire \cmd_mux|src_data[35]~combout ;
wire \cmd_mux|src_data[34]~combout ;
wire \cmd_mux|src_data[33]~combout ;
wire \cmd_mux|src_data[32]~combout ;
wire \link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ;
wire \link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ;
wire \link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ;
wire \link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ;
wire \link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ;
wire \link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ;
wire \flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ;
wire \router_001|Equal4~0_combout ;
wire \hps_0_h2f_axi_master_rd_limiter|last_channel[4]~q ;
wire \cmd_mux_004|src_valid~0_combout ;
wire \flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ;
wire \flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ;
wire \flags_s1_agent_rsp_fifo|write~0_combout ;
wire \flags_s1_agent_rsp_fifo|write~1_combout ;
wire \tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ;
wire \router_001|Equal7~0_combout ;
wire \hps_0_h2f_axi_master_rd_limiter|last_channel[7]~q ;
wire \cmd_mux_007|src_valid~0_combout ;
wire \tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ;
wire \tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ;
wire \tx_full_s1_agent_rsp_fifo|write~0_combout ;
wire \tx_full_s1_agent_rsp_fifo|write~1_combout ;
wire \flags_s1_agent|cp_ready~1_combout ;
wire \flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ;
wire \flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ;
wire \flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ;
wire \flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ;
wire \flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ;
wire \tx_full_s1_agent|cp_ready~1_combout ;
wire \tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ;
wire \tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ;
wire \tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ;
wire \tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ;
wire \tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ;
wire \autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ;
wire \hps_0_h2f_axi_master_wr_limiter|last_channel[2]~q ;
wire \cmd_demux|src2_valid~0_combout ;
wire \cmd_demux|src2_valid~1_combout ;
wire \router_001|src_channel[2]~4_combout ;
wire \hps_0_h2f_axi_master_rd_limiter|last_channel[2]~q ;
wire \cmd_demux_001|src2_valid~0_combout ;
wire \cmd_mux_002|src_valid~0_combout ;
wire \autostart_s1_agent|cp_ready~3_combout ;
wire \autostart_s1_agent|uncompressor|last_packet_beat~2_combout ;
wire \rsp_demux_002|WideOr0~0_combout ;
wire \autostart_s1_agent_rsp_fifo|read~0_combout ;
wire \autostart_s1_agent|cp_ready~4_combout ;
wire \autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ;
wire \autostart_s1_agent|rf_source_valid~0_combout ;
wire \cmd_mux_002|src_data[87]~combout ;
wire \cmd_mux_002|src_data[88]~combout ;
wire \cmd_mux_002|src_valid~1_combout ;
wire \cmd_mux_002|src_data[35]~combout ;
wire \cmd_mux_002|src_data[34]~combout ;
wire \cmd_mux_002|src_data[33]~combout ;
wire \cmd_mux_002|src_data[32]~combout ;
wire \autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ;
wire \autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ;
wire \autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ;
wire \autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ;
wire \autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ;
wire \autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ;
wire \cmd_mux_002|src_payload[0]~combout ;
wire \cmd_demux|src2_valid~2_combout ;
wire \cmd_demux_001|src2_valid~1_combout ;
wire \wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ;
wire \cmd_demux|src6_valid~0_combout ;
wire \cmd_demux|src6_valid~1_combout ;
wire \cmd_demux_001|src6_valid~0_combout ;
wire \cmd_mux_006|src_valid~0_combout ;
wire \wr_data_s1_agent|cp_ready~3_combout ;
wire \wr_data_s1_agent|uncompressor|last_packet_beat~2_combout ;
wire \rsp_demux_006|WideOr0~0_combout ;
wire \wr_data_s1_agent_rsp_fifo|read~0_combout ;
wire \wr_data_s1_agent|cp_ready~4_combout ;
wire \wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ;
wire \wr_data_s1_agent|rf_source_valid~0_combout ;
wire \cmd_mux_006|src_data[87]~combout ;
wire \cmd_mux_006|src_data[88]~combout ;
wire \cmd_mux_006|src_valid~1_combout ;
wire \cmd_mux_006|src_data[35]~combout ;
wire \cmd_mux_006|src_data[34]~combout ;
wire \cmd_mux_006|src_data[33]~combout ;
wire \cmd_mux_006|src_data[32]~combout ;
wire \wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ;
wire \wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ;
wire \wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ;
wire \wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ;
wire \wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ;
wire \wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ;
wire \cmd_mux_006|src_payload[0]~combout ;
wire \cmd_demux|src6_valid~2_combout ;
wire \cmd_demux_001|src6_valid~1_combout ;
wire \rsp_mux|src_payload~0_combout ;
wire \rsp_mux|src_payload~1_combout ;
wire \rsp_mux|src_payload[0]~8_combout ;
wire \rsp_mux|src_payload[0]~9_combout ;
wire \router|Equal6~0_combout ;
wire \wr_data_s1_agent|uncompressor|sink_ready~0_combout ;
wire \rd_data_s1_agent|uncompressor|sink_ready~0_combout ;
wire \link_start_s1_agent|uncompressor|sink_ready~0_combout ;
wire \link_disable_s1_agent|uncompressor|sink_ready~0_combout ;
wire \autostart_s1_agent|uncompressor|sink_ready~0_combout ;
wire \data_i_s1_agent|uncompressor|sink_ready~0_combout ;
wire \tick_in_s1_agent|rp_valid~combout ;
wire \time_in_s1_agent|rp_valid~combout ;
wire \tx_clk_div_s1_agent|uncompressor|sink_ready~0_combout ;
wire \spill_enable_s1_agent|uncompressor|sink_ready~0_combout ;
wire \tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ;
wire \spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ;
wire \tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ;
wire \time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ;
wire \autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ;
wire \rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ;
wire \link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ;
wire \link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ;
wire \data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ;
wire \wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ;
wire \tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ;
wire \spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ;
wire \tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ;
wire \time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ;
wire \autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ;
wire \rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ;
wire \link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ;
wire \link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ;
wire \data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ;
wire \wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ;
wire \tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ;
wire \spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ;
wire \tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ;
wire \time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ;
wire \autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ;
wire \rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ;
wire \link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ;
wire \link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ;
wire \data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ;
wire \wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ;
wire \tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ;
wire \spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ;
wire \tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ;
wire \time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ;
wire \autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ;
wire \rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ;
wire \link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ;
wire \link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ;
wire \data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ;
wire \wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ;
wire \tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ;
wire \spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ;
wire \tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ;
wire \time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ;
wire \autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ;
wire \rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ;
wire \link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ;
wire \link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ;
wire \data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ;
wire \wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ;
wire \tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ;
wire \spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ;
wire \tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ;
wire \time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ;
wire \autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ;
wire \rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ;
wire \link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ;
wire \link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ;
wire \data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ;
wire \wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ;
wire \tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ;
wire \spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ;
wire \tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ;
wire \time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ;
wire \autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ;
wire \rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ;
wire \link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ;
wire \link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ;
wire \data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ;
wire \wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ;
wire \tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ;
wire \spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ;
wire \tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ;
wire \time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ;
wire \autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ;
wire \rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ;
wire \link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ;
wire \link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ;
wire \data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ;
wire \wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ;
wire \tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ;
wire \spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ;
wire \tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ;
wire \time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ;
wire \autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ;
wire \rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ;
wire \link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ;
wire \link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ;
wire \data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ;
wire \wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ;
wire \tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ;
wire \spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ;
wire \tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ;
wire \time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ;
wire \autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ;
wire \rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ;
wire \link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ;
wire \link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ;
wire \data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ;
wire \wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ;
wire \tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ;
wire \spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ;
wire \tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ;
wire \time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ;
wire \autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ;
wire \rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ;
wire \link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ;
wire \link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ;
wire \data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ;
wire \wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ;
wire \tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ;
wire \spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ;
wire \tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ;
wire \time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ;
wire \autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ;
wire \rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ;
wire \link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ;
wire \link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ;
wire \data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ;
wire \wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ;
wire \time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ;
wire \currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ;
wire \flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ;
wire \tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ;
wire \data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ;
wire \rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ;
wire \tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ;
wire \time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ;
wire \currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ;
wire \flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ;
wire \tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ;
wire \data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ;
wire \rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ;
wire \tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ;
wire \time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ;
wire \currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ;
wire \flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ;
wire \tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ;
wire \data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ;
wire \rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ;
wire \tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ;
wire \time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ;
wire \currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ;
wire \flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ;
wire \tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ;
wire \data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ;
wire \rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ;
wire \tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ;
wire \time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ;
wire \currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ;
wire \flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ;
wire \tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ;
wire \data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ;
wire \rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ;
wire \tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ;
wire \time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ;
wire \currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ;
wire \flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ;
wire \tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ;
wire \data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ;
wire \rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ;
wire \tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ;
wire \time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ;
wire \currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ;
wire \flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ;
wire \tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ;
wire \data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ;
wire \rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ;
wire \tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ;
wire \time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ;
wire \currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ;
wire \flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ;
wire \tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ;
wire \data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ;
wire \rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ;
wire \tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ;
wire \time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ;
wire \currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ;
wire \flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ;
wire \tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ;
wire \data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ;
wire \rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ;
wire \tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ;
wire \time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ;
wire \currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ;
wire \flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ;
wire \tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ;
wire \data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ;
wire \rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ;
wire \tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ;
wire \time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ;
wire \currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ;
wire \flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ;
wire \tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ;
wire \data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ;
wire \rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ;
wire \tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ;
wire \time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ;
wire \currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ;
wire \flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ;
wire \tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ;
wire \data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ;
wire \rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ;
wire \tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ;
wire \cmd_mux_002|src_payload~0_combout ;
wire \hps_0_h2f_axi_master_agent|Selector3~0_combout ;
wire \hps_0_h2f_axi_master_agent|Selector10~0_combout ;
wire \hps_0_h2f_axi_master_agent|Selector10~1_combout ;
wire \cmd_mux_002|src_data[82]~combout ;
wire \hps_0_h2f_axi_master_agent|align_address_to_size|base_address[3]~0_combout ;
wire \hps_0_h2f_axi_master_agent|Selector4~1_combout ;
wire \hps_0_h2f_axi_master_agent|Add3~1_combout ;
wire \hps_0_h2f_axi_master_agent|Add3~2_combout ;
wire \hps_0_h2f_axi_master_agent|Selector11~0_combout ;
wire \hps_0_h2f_axi_master_agent|Selector11~1_combout ;
wire \cmd_mux_002|src_data[81]~combout ;
wire \hps_0_h2f_axi_master_agent|align_address_to_size|base_address[2]~1_combout ;
wire \cmd_mux_005|src_payload~0_combout ;
wire \cmd_mux_005|src_data[82]~combout ;
wire \cmd_mux_005|src_data[81]~combout ;
wire \cmd_mux_005|src_payload~1_combout ;
wire \cmd_mux_005|src_payload~2_combout ;
wire \cmd_mux_005|src_payload~3_combout ;
wire \cmd_mux_005|src_payload~4_combout ;
wire \cmd_mux_005|src_payload~5_combout ;
wire \cmd_mux_005|src_payload~6_combout ;
wire \cmd_mux_005|src_payload~7_combout ;
wire \cmd_mux_005|src_payload~8_combout ;
wire \cmd_mux_001|src_payload~0_combout ;
wire \cmd_mux_001|src_data[82]~combout ;
wire \cmd_mux_001|src_data[81]~combout ;
wire \cmd_mux|src_payload~0_combout ;
wire \cmd_mux|src_data[82]~combout ;
wire \cmd_mux|src_data[81]~combout ;
wire \cmd_mux_009|src_payload~0_combout ;
wire \cmd_mux_009|src_data[82]~combout ;
wire \cmd_mux_009|src_data[81]~combout ;
wire \cmd_mux_016|src_payload~0_combout ;
wire \cmd_mux_016|src_data[82]~combout ;
wire \cmd_mux_016|src_data[81]~combout ;
wire \cmd_mux_013|src_payload~0_combout ;
wire \cmd_mux_013|src_data[82]~combout ;
wire \cmd_mux_013|src_data[81]~combout ;
wire \cmd_mux_014|src_payload~0_combout ;
wire \cmd_mux_014|src_data[82]~combout ;
wire \cmd_mux_014|src_data[81]~combout ;
wire \cmd_mux_014|src_payload~1_combout ;
wire \cmd_mux_014|src_payload~2_combout ;
wire \cmd_mux_014|src_payload~3_combout ;
wire \cmd_mux_014|src_payload~4_combout ;
wire \cmd_mux_014|src_payload~5_combout ;
wire \cmd_mux_014|src_payload~6_combout ;
wire \cmd_mux_014|src_payload~7_combout ;
wire \cmd_mux_015|src_payload~0_combout ;
wire \cmd_mux_015|src_data[82]~combout ;
wire \cmd_mux_015|src_data[81]~combout ;
wire \cmd_mux_015|src_payload~1_combout ;
wire \cmd_mux_015|src_payload~2_combout ;
wire \cmd_mux_015|src_payload~3_combout ;
wire \cmd_mux_015|src_payload~4_combout ;
wire \cmd_mux_015|src_payload~5_combout ;
wire \cmd_mux_015|src_payload~6_combout ;
wire \cmd_mux_006|src_payload~0_combout ;
wire \cmd_mux_006|src_data[82]~combout ;
wire \cmd_mux_006|src_data[81]~combout ;
wire \router|src_channel~0_combout ;
wire \router|Equal15~2_combout ;
wire \router|Equal16~2_combout ;
wire \router|Equal13~1_combout ;
wire \router|Equal14~2_combout ;
wire \router|Equal5~2_combout ;
wire \router_001|src_channel~5_combout ;
wire \router|Equal9~1_combout ;
wire \router|src_channel[0]~1_combout ;
wire \router|Equal2~0_combout ;
wire \cmd_mux_015|src_data[105]~combout ;
wire \cmd_mux_016|src_data[105]~combout ;
wire \cmd_mux_013|src_data[105]~combout ;
wire \cmd_mux_014|src_data[105]~combout ;
wire \cmd_mux_002|src_data[105]~combout ;
wire \cmd_mux_009|src_data[105]~combout ;
wire \cmd_mux|src_data[105]~combout ;
wire \cmd_mux_001|src_data[105]~combout ;
wire \cmd_mux_005|src_data[105]~combout ;
wire \cmd_mux_006|src_data[105]~combout ;
wire \cmd_mux_015|src_data[106]~combout ;
wire \cmd_mux_016|src_data[106]~combout ;
wire \cmd_mux_013|src_data[106]~combout ;
wire \cmd_mux_014|src_data[106]~combout ;
wire \cmd_mux_002|src_data[106]~combout ;
wire \cmd_mux_009|src_data[106]~combout ;
wire \cmd_mux|src_data[106]~combout ;
wire \cmd_mux_001|src_data[106]~combout ;
wire \cmd_mux_005|src_data[106]~combout ;
wire \cmd_mux_006|src_data[106]~combout ;
wire \cmd_mux_015|src_data[107]~combout ;
wire \cmd_mux_016|src_data[107]~combout ;
wire \cmd_mux_013|src_data[107]~combout ;
wire \cmd_mux_014|src_data[107]~combout ;
wire \cmd_mux_002|src_data[107]~combout ;
wire \cmd_mux_009|src_data[107]~combout ;
wire \cmd_mux|src_data[107]~combout ;
wire \cmd_mux_001|src_data[107]~combout ;
wire \cmd_mux_005|src_data[107]~combout ;
wire \cmd_mux_006|src_data[107]~combout ;
wire \cmd_mux_015|src_data[108]~combout ;
wire \cmd_mux_016|src_data[108]~combout ;
wire \cmd_mux_013|src_data[108]~combout ;
wire \cmd_mux_014|src_data[108]~combout ;
wire \cmd_mux_002|src_data[108]~combout ;
wire \cmd_mux_009|src_data[108]~combout ;
wire \cmd_mux|src_data[108]~combout ;
wire \cmd_mux_001|src_data[108]~combout ;
wire \cmd_mux_005|src_data[108]~combout ;
wire \cmd_mux_006|src_data[108]~combout ;
wire \cmd_mux_015|src_data[109]~combout ;
wire \cmd_mux_016|src_data[109]~combout ;
wire \cmd_mux_013|src_data[109]~combout ;
wire \cmd_mux_014|src_data[109]~combout ;
wire \cmd_mux_002|src_data[109]~combout ;
wire \cmd_mux_009|src_data[109]~combout ;
wire \cmd_mux|src_data[109]~combout ;
wire \cmd_mux_001|src_data[109]~combout ;
wire \cmd_mux_005|src_data[109]~combout ;
wire \cmd_mux_006|src_data[109]~combout ;
wire \cmd_mux_015|src_data[110]~combout ;
wire \cmd_mux_016|src_data[110]~combout ;
wire \cmd_mux_013|src_data[110]~combout ;
wire \cmd_mux_014|src_data[110]~combout ;
wire \cmd_mux_002|src_data[110]~combout ;
wire \cmd_mux_009|src_data[110]~combout ;
wire \cmd_mux|src_data[110]~combout ;
wire \cmd_mux_001|src_data[110]~combout ;
wire \cmd_mux_005|src_data[110]~combout ;
wire \cmd_mux_006|src_data[110]~combout ;
wire \cmd_mux_015|src_data[111]~combout ;
wire \cmd_mux_016|src_data[111]~combout ;
wire \cmd_mux_013|src_data[111]~combout ;
wire \cmd_mux_014|src_data[111]~combout ;
wire \cmd_mux_002|src_data[111]~combout ;
wire \cmd_mux_009|src_data[111]~combout ;
wire \cmd_mux|src_data[111]~combout ;
wire \cmd_mux_001|src_data[111]~combout ;
wire \cmd_mux_005|src_data[111]~combout ;
wire \cmd_mux_006|src_data[111]~combout ;
wire \cmd_mux_015|src_data[112]~combout ;
wire \cmd_mux_016|src_data[112]~combout ;
wire \cmd_mux_013|src_data[112]~combout ;
wire \cmd_mux_014|src_data[112]~combout ;
wire \cmd_mux_002|src_data[112]~combout ;
wire \cmd_mux_009|src_data[112]~combout ;
wire \cmd_mux|src_data[112]~combout ;
wire \cmd_mux_001|src_data[112]~combout ;
wire \cmd_mux_005|src_data[112]~combout ;
wire \cmd_mux_006|src_data[112]~combout ;
wire \cmd_mux_015|src_data[113]~combout ;
wire \cmd_mux_016|src_data[113]~combout ;
wire \cmd_mux_013|src_data[113]~combout ;
wire \cmd_mux_014|src_data[113]~combout ;
wire \cmd_mux_002|src_data[113]~combout ;
wire \cmd_mux_009|src_data[113]~combout ;
wire \cmd_mux|src_data[113]~combout ;
wire \cmd_mux_001|src_data[113]~combout ;
wire \cmd_mux_005|src_data[113]~combout ;
wire \cmd_mux_006|src_data[113]~combout ;
wire \cmd_mux_015|src_data[114]~combout ;
wire \cmd_mux_016|src_data[114]~combout ;
wire \cmd_mux_013|src_data[114]~combout ;
wire \cmd_mux_014|src_data[114]~combout ;
wire \cmd_mux_002|src_data[114]~combout ;
wire \cmd_mux_009|src_data[114]~combout ;
wire \cmd_mux|src_data[114]~combout ;
wire \cmd_mux_001|src_data[114]~combout ;
wire \cmd_mux_005|src_data[114]~combout ;
wire \cmd_mux_006|src_data[114]~combout ;
wire \cmd_mux_015|src_data[115]~combout ;
wire \cmd_mux_016|src_data[115]~combout ;
wire \cmd_mux_013|src_data[115]~combout ;
wire \cmd_mux_014|src_data[115]~combout ;
wire \cmd_mux_002|src_data[115]~combout ;
wire \cmd_mux_009|src_data[115]~combout ;
wire \cmd_mux|src_data[115]~combout ;
wire \cmd_mux_001|src_data[115]~combout ;
wire \cmd_mux_005|src_data[115]~combout ;
wire \cmd_mux_006|src_data[115]~combout ;
wire \cmd_mux_015|src_data[116]~combout ;
wire \cmd_mux_016|src_data[116]~combout ;
wire \cmd_mux_013|src_data[116]~combout ;
wire \cmd_mux_014|src_data[116]~combout ;
wire \cmd_mux_002|src_data[116]~combout ;
wire \cmd_mux_009|src_data[116]~combout ;
wire \cmd_mux|src_data[116]~combout ;
wire \cmd_mux_001|src_data[116]~combout ;
wire \cmd_mux_005|src_data[116]~combout ;
wire \cmd_mux_006|src_data[116]~combout ;
wire \cmd_mux_002|src_data[86]~combout ;
wire \cmd_mux_005|src_data[86]~combout ;
wire \cmd_mux_001|src_data[86]~combout ;
wire \cmd_mux|src_data[86]~combout ;
wire \cmd_mux_009|src_data[86]~combout ;
wire \cmd_mux_016|src_data[86]~combout ;
wire \cmd_mux_013|src_data[86]~combout ;
wire \cmd_mux_014|src_data[86]~combout ;
wire \cmd_mux_015|src_data[86]~combout ;
wire \cmd_mux_006|src_data[86]~combout ;
wire \hps_0_h2f_axi_master_agent|Selector5~1_combout ;
wire \hps_0_h2f_axi_master_agent|Add3~3_combout ;
wire \hps_0_h2f_axi_master_agent|Selector12~0_combout ;
wire \cmd_mux_002|src_data[80]~combout ;
wire \hps_0_h2f_axi_master_agent|align_address_to_size|out_data[1]~5_combout ;
wire \cmd_mux_005|src_data[80]~combout ;
wire \cmd_mux_001|src_data[80]~combout ;
wire \cmd_mux|src_data[80]~combout ;
wire \cmd_mux_009|src_data[80]~combout ;
wire \cmd_mux_016|src_data[80]~combout ;
wire \cmd_mux_013|src_data[80]~combout ;
wire \cmd_mux_014|src_data[80]~combout ;
wire \cmd_mux_015|src_data[80]~combout ;
wire \cmd_mux_006|src_data[80]~combout ;
wire \cmd_mux_003|src_payload~0_combout ;
wire \cmd_mux_003|src_payload~1_combout ;
wire \cmd_mux_003|src_payload~2_combout ;
wire \cmd_mux_008|src_payload~0_combout ;
wire \cmd_mux_008|src_payload~1_combout ;
wire \cmd_mux_008|src_payload~2_combout ;
wire \cmd_mux_007|src_payload~0_combout ;
wire \cmd_mux_007|src_payload~1_combout ;
wire \cmd_mux_007|src_payload~2_combout ;
wire \cmd_mux_004|src_payload~0_combout ;
wire \cmd_mux_004|src_payload~1_combout ;
wire \cmd_mux_004|src_payload~2_combout ;
wire \cmd_mux_012|src_payload~0_combout ;
wire \cmd_mux_012|src_payload~1_combout ;
wire \cmd_mux_012|src_payload~2_combout ;
wire \cmd_mux_011|src_payload~0_combout ;
wire \cmd_mux_011|src_payload~1_combout ;
wire \cmd_mux_011|src_payload~2_combout ;
wire \cmd_mux_010|src_payload~0_combout ;
wire \cmd_mux_010|src_payload~1_combout ;
wire \cmd_mux_010|src_payload~2_combout ;
wire \hps_0_h2f_axi_master_agent|align_address_to_size|out_data[0]~6_combout ;
wire \hps_0_h2f_axi_master_agent|Selector6~0_combout ;
wire \hps_0_h2f_axi_master_agent|Selector13~1_combout ;
wire \cmd_mux_002|src_data[79]~combout ;
wire \cmd_mux_005|src_data[79]~combout ;
wire \cmd_mux_001|src_data[79]~combout ;
wire \cmd_mux|src_data[79]~combout ;
wire \cmd_mux_009|src_data[79]~combout ;
wire \cmd_mux_016|src_data[79]~combout ;
wire \cmd_mux_013|src_data[79]~combout ;
wire \cmd_mux_014|src_data[79]~combout ;
wire \cmd_mux_015|src_data[79]~combout ;
wire \cmd_mux_006|src_data[79]~combout ;
wire \time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_burstwrap[1]~0_combout ;
wire \time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_addr[2]~2_combout ;


spw_babasu_spw_babasu_mm_interconnect_0_cmd_mux_9 cmd_mux_009(
	.h2f_WLAST_0(h2f_WLAST_0),
	.h2f_ARID_0(h2f_ARID_0),
	.h2f_ARID_1(h2f_ARID_1),
	.h2f_ARID_2(h2f_ARID_2),
	.h2f_ARID_3(h2f_ARID_3),
	.h2f_ARID_4(h2f_ARID_4),
	.h2f_ARID_5(h2f_ARID_5),
	.h2f_ARID_6(h2f_ARID_6),
	.h2f_ARID_7(h2f_ARID_7),
	.h2f_ARID_8(h2f_ARID_8),
	.h2f_ARID_9(h2f_ARID_9),
	.h2f_ARID_10(h2f_ARID_10),
	.h2f_ARID_11(h2f_ARID_11),
	.h2f_ARSIZE_0(h2f_ARSIZE_0),
	.h2f_ARSIZE_1(h2f_ARSIZE_1),
	.h2f_ARSIZE_2(h2f_ARSIZE_2),
	.h2f_AWID_0(h2f_AWID_0),
	.h2f_AWID_1(h2f_AWID_1),
	.h2f_AWID_2(h2f_AWID_2),
	.h2f_AWID_3(h2f_AWID_3),
	.h2f_AWID_4(h2f_AWID_4),
	.h2f_AWID_5(h2f_AWID_5),
	.h2f_AWID_6(h2f_AWID_6),
	.h2f_AWID_7(h2f_AWID_7),
	.h2f_AWID_8(h2f_AWID_8),
	.h2f_AWID_9(h2f_AWID_9),
	.h2f_AWID_10(h2f_AWID_10),
	.h2f_AWID_11(h2f_AWID_11),
	.h2f_AWSIZE_0(h2f_AWSIZE_0),
	.h2f_AWSIZE_1(h2f_AWSIZE_1),
	.h2f_AWSIZE_2(h2f_AWSIZE_2),
	.h2f_WDATA_0(h2f_WDATA_0),
	.h2f_WSTRB_0(h2f_WSTRB_0),
	.h2f_WSTRB_1(h2f_WSTRB_1),
	.h2f_WSTRB_2(h2f_WSTRB_2),
	.h2f_WSTRB_3(h2f_WSTRB_3),
	.nxt_in_ready(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.nxt_in_ready1(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.saved_grant_1(\cmd_mux_009|saved_grant[1]~q ),
	.write_addr_data_both_valid(\hps_0_h2f_axi_master_agent|write_addr_data_both_valid~combout ),
	.out_data_5(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[5]~1_combout ),
	.Equal15(\router|Equal15~0_combout ),
	.Equal9(\router|Equal9~0_combout ),
	.saved_grant_0(\cmd_mux_009|saved_grant[0]~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.Equal5(\router|Equal5~1_combout ),
	.src9_valid(\cmd_demux|src9_valid~0_combout ),
	.src9_valid1(\cmd_demux|src9_valid~1_combout ),
	.Equal91(\router_001|Equal9~0_combout ),
	.src9_valid2(\cmd_demux_001|src9_valid~0_combout ),
	.src_valid(\cmd_mux_009|src_valid~0_combout ),
	.src_data_87(\cmd_mux_009|src_data[87]~combout ),
	.src_data_88(\cmd_mux_009|src_data[88]~combout ),
	.src_valid1(\cmd_mux_009|src_valid~1_combout ),
	.src_data_35(\cmd_mux_009|src_data[35]~combout ),
	.src_data_34(\cmd_mux_009|src_data[34]~combout ),
	.src_data_33(\cmd_mux_009|src_data[33]~combout ),
	.src_data_32(\cmd_mux_009|src_data[32]~combout ),
	.src_payload_0(\cmd_mux_009|src_payload[0]~combout ),
	.src9_valid3(\cmd_demux|src9_valid~2_combout ),
	.src9_valid4(\cmd_demux_001|src9_valid~1_combout ),
	.Selector3(\hps_0_h2f_axi_master_agent|Selector3~0_combout ),
	.Selector10(\hps_0_h2f_axi_master_agent|Selector10~1_combout ),
	.Selector4(\hps_0_h2f_axi_master_agent|Selector4~1_combout ),
	.Selector11(\hps_0_h2f_axi_master_agent|Selector11~1_combout ),
	.src_payload(\cmd_mux_009|src_payload~0_combout ),
	.src_data_82(\cmd_mux_009|src_data[82]~combout ),
	.src_data_81(\cmd_mux_009|src_data[81]~combout ),
	.src_data_105(\cmd_mux_009|src_data[105]~combout ),
	.src_data_106(\cmd_mux_009|src_data[106]~combout ),
	.src_data_107(\cmd_mux_009|src_data[107]~combout ),
	.src_data_108(\cmd_mux_009|src_data[108]~combout ),
	.src_data_109(\cmd_mux_009|src_data[109]~combout ),
	.src_data_110(\cmd_mux_009|src_data[110]~combout ),
	.src_data_111(\cmd_mux_009|src_data[111]~combout ),
	.src_data_112(\cmd_mux_009|src_data[112]~combout ),
	.src_data_113(\cmd_mux_009|src_data[113]~combout ),
	.src_data_114(\cmd_mux_009|src_data[114]~combout ),
	.src_data_115(\cmd_mux_009|src_data[115]~combout ),
	.src_data_116(\cmd_mux_009|src_data[116]~combout ),
	.src_data_86(\cmd_mux_009|src_data[86]~combout ),
	.Selector5(\hps_0_h2f_axi_master_agent|Selector5~1_combout ),
	.Selector12(\hps_0_h2f_axi_master_agent|Selector12~0_combout ),
	.src_data_80(\cmd_mux_009|src_data[80]~combout ),
	.Selector6(\hps_0_h2f_axi_master_agent|Selector6~0_combout ),
	.Selector13(\hps_0_h2f_axi_master_agent|Selector13~1_combout ),
	.src_data_79(\cmd_mux_009|src_data[79]~combout ),
	.clk_clk(clk_clk));

spw_babasu_spw_babasu_mm_interconnect_0_cmd_mux_8 cmd_mux_008(
	.h2f_ARVALID_0(h2f_ARVALID_0),
	.h2f_ARSIZE_0(h2f_ARSIZE_0),
	.h2f_ARSIZE_1(h2f_ARSIZE_1),
	.h2f_ARSIZE_2(h2f_ARSIZE_2),
	.has_pending_responses(\hps_0_h2f_axi_master_rd_limiter|has_pending_responses~q ),
	.saved_grant_1(\cmd_mux_008|saved_grant[1]~q ),
	.src_channel(\router_001|src_channel~0_combout ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.nxt_in_ready(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.last_channel_8(\hps_0_h2f_axi_master_rd_limiter|last_channel[8]~q ),
	.src_valid(\cmd_mux_008|src_valid~0_combout ),
	.src_payload(\cmd_mux_008|src_payload~0_combout ),
	.src_payload1(\cmd_mux_008|src_payload~1_combout ),
	.src_payload2(\cmd_mux_008|src_payload~2_combout ),
	.clk_clk(clk_clk));

spw_babasu_spw_babasu_mm_interconnect_0_cmd_mux_7 cmd_mux_007(
	.h2f_ARVALID_0(h2f_ARVALID_0),
	.h2f_ARSIZE_0(h2f_ARSIZE_0),
	.h2f_ARSIZE_1(h2f_ARSIZE_1),
	.h2f_ARSIZE_2(h2f_ARSIZE_2),
	.has_pending_responses(\hps_0_h2f_axi_master_rd_limiter|has_pending_responses~q ),
	.saved_grant_1(\cmd_mux_007|saved_grant[1]~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.nxt_in_ready(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ),
	.Equal7(\router_001|Equal7~0_combout ),
	.last_channel_7(\hps_0_h2f_axi_master_rd_limiter|last_channel[7]~q ),
	.src_valid(\cmd_mux_007|src_valid~0_combout ),
	.src_payload(\cmd_mux_007|src_payload~0_combout ),
	.src_payload1(\cmd_mux_007|src_payload~1_combout ),
	.src_payload2(\cmd_mux_007|src_payload~2_combout ),
	.clk_clk(clk_clk));

spw_babasu_spw_babasu_mm_interconnect_0_cmd_mux_6 cmd_mux_006(
	.h2f_WLAST_0(h2f_WLAST_0),
	.h2f_ARID_0(h2f_ARID_0),
	.h2f_ARID_1(h2f_ARID_1),
	.h2f_ARID_2(h2f_ARID_2),
	.h2f_ARID_3(h2f_ARID_3),
	.h2f_ARID_4(h2f_ARID_4),
	.h2f_ARID_5(h2f_ARID_5),
	.h2f_ARID_6(h2f_ARID_6),
	.h2f_ARID_7(h2f_ARID_7),
	.h2f_ARID_8(h2f_ARID_8),
	.h2f_ARID_9(h2f_ARID_9),
	.h2f_ARID_10(h2f_ARID_10),
	.h2f_ARID_11(h2f_ARID_11),
	.h2f_ARSIZE_0(h2f_ARSIZE_0),
	.h2f_ARSIZE_1(h2f_ARSIZE_1),
	.h2f_ARSIZE_2(h2f_ARSIZE_2),
	.h2f_AWID_0(h2f_AWID_0),
	.h2f_AWID_1(h2f_AWID_1),
	.h2f_AWID_2(h2f_AWID_2),
	.h2f_AWID_3(h2f_AWID_3),
	.h2f_AWID_4(h2f_AWID_4),
	.h2f_AWID_5(h2f_AWID_5),
	.h2f_AWID_6(h2f_AWID_6),
	.h2f_AWID_7(h2f_AWID_7),
	.h2f_AWID_8(h2f_AWID_8),
	.h2f_AWID_9(h2f_AWID_9),
	.h2f_AWID_10(h2f_AWID_10),
	.h2f_AWID_11(h2f_AWID_11),
	.h2f_AWSIZE_0(h2f_AWSIZE_0),
	.h2f_AWSIZE_1(h2f_AWSIZE_1),
	.h2f_AWSIZE_2(h2f_AWSIZE_2),
	.h2f_WDATA_0(h2f_WDATA_0),
	.h2f_WSTRB_0(h2f_WSTRB_0),
	.h2f_WSTRB_1(h2f_WSTRB_1),
	.h2f_WSTRB_2(h2f_WSTRB_2),
	.h2f_WSTRB_3(h2f_WSTRB_3),
	.nxt_in_ready(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.Equal6(\router_001|Equal6~0_combout ),
	.nxt_in_ready1(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.saved_grant_1(\cmd_mux_006|saved_grant[1]~q ),
	.write_addr_data_both_valid(\hps_0_h2f_axi_master_agent|write_addr_data_both_valid~combout ),
	.out_data_4(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[4]~2_combout ),
	.Equal5(\router|Equal5~0_combout ),
	.Equal14(\router|Equal14~0_combout ),
	.saved_grant_0(\cmd_mux_006|saved_grant[0]~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.Equal141(\router|Equal14~1_combout ),
	.src6_valid(\cmd_demux|src6_valid~0_combout ),
	.src6_valid1(\cmd_demux|src6_valid~1_combout ),
	.src6_valid2(\cmd_demux_001|src6_valid~0_combout ),
	.src_valid(\cmd_mux_006|src_valid~0_combout ),
	.src_data_87(\cmd_mux_006|src_data[87]~combout ),
	.src_data_88(\cmd_mux_006|src_data[88]~combout ),
	.src_valid1(\cmd_mux_006|src_valid~1_combout ),
	.src_data_35(\cmd_mux_006|src_data[35]~combout ),
	.src_data_34(\cmd_mux_006|src_data[34]~combout ),
	.src_data_33(\cmd_mux_006|src_data[33]~combout ),
	.src_data_32(\cmd_mux_006|src_data[32]~combout ),
	.src_payload_0(\cmd_mux_006|src_payload[0]~combout ),
	.src6_valid3(\cmd_demux|src6_valid~2_combout ),
	.src6_valid4(\cmd_demux_001|src6_valid~1_combout ),
	.Selector3(\hps_0_h2f_axi_master_agent|Selector3~0_combout ),
	.Selector10(\hps_0_h2f_axi_master_agent|Selector10~1_combout ),
	.Selector4(\hps_0_h2f_axi_master_agent|Selector4~1_combout ),
	.Selector11(\hps_0_h2f_axi_master_agent|Selector11~1_combout ),
	.src_payload(\cmd_mux_006|src_payload~0_combout ),
	.src_data_82(\cmd_mux_006|src_data[82]~combout ),
	.src_data_81(\cmd_mux_006|src_data[81]~combout ),
	.src_data_105(\cmd_mux_006|src_data[105]~combout ),
	.src_data_106(\cmd_mux_006|src_data[106]~combout ),
	.src_data_107(\cmd_mux_006|src_data[107]~combout ),
	.src_data_108(\cmd_mux_006|src_data[108]~combout ),
	.src_data_109(\cmd_mux_006|src_data[109]~combout ),
	.src_data_110(\cmd_mux_006|src_data[110]~combout ),
	.src_data_111(\cmd_mux_006|src_data[111]~combout ),
	.src_data_112(\cmd_mux_006|src_data[112]~combout ),
	.src_data_113(\cmd_mux_006|src_data[113]~combout ),
	.src_data_114(\cmd_mux_006|src_data[114]~combout ),
	.src_data_115(\cmd_mux_006|src_data[115]~combout ),
	.src_data_116(\cmd_mux_006|src_data[116]~combout ),
	.src_data_86(\cmd_mux_006|src_data[86]~combout ),
	.Selector5(\hps_0_h2f_axi_master_agent|Selector5~1_combout ),
	.Selector12(\hps_0_h2f_axi_master_agent|Selector12~0_combout ),
	.src_data_80(\cmd_mux_006|src_data[80]~combout ),
	.Selector6(\hps_0_h2f_axi_master_agent|Selector6~0_combout ),
	.Selector13(\hps_0_h2f_axi_master_agent|Selector13~1_combout ),
	.src_data_79(\cmd_mux_006|src_data[79]~combout ),
	.clk_clk(clk_clk));

spw_babasu_spw_babasu_mm_interconnect_0_cmd_mux_5 cmd_mux_005(
	.h2f_ARVALID_0(h2f_ARVALID_0),
	.h2f_WLAST_0(h2f_WLAST_0),
	.h2f_ARADDR_4(h2f_ARADDR_4),
	.h2f_ARADDR_5(h2f_ARADDR_5),
	.h2f_ARADDR_6(h2f_ARADDR_6),
	.h2f_ARADDR_7(h2f_ARADDR_7),
	.h2f_ARADDR_8(h2f_ARADDR_8),
	.h2f_ARID_0(h2f_ARID_0),
	.h2f_ARID_1(h2f_ARID_1),
	.h2f_ARID_2(h2f_ARID_2),
	.h2f_ARID_3(h2f_ARID_3),
	.h2f_ARID_4(h2f_ARID_4),
	.h2f_ARID_5(h2f_ARID_5),
	.h2f_ARID_6(h2f_ARID_6),
	.h2f_ARID_7(h2f_ARID_7),
	.h2f_ARID_8(h2f_ARID_8),
	.h2f_ARID_9(h2f_ARID_9),
	.h2f_ARID_10(h2f_ARID_10),
	.h2f_ARID_11(h2f_ARID_11),
	.h2f_ARSIZE_0(h2f_ARSIZE_0),
	.h2f_ARSIZE_1(h2f_ARSIZE_1),
	.h2f_ARSIZE_2(h2f_ARSIZE_2),
	.h2f_AWID_0(h2f_AWID_0),
	.h2f_AWID_1(h2f_AWID_1),
	.h2f_AWID_2(h2f_AWID_2),
	.h2f_AWID_3(h2f_AWID_3),
	.h2f_AWID_4(h2f_AWID_4),
	.h2f_AWID_5(h2f_AWID_5),
	.h2f_AWID_6(h2f_AWID_6),
	.h2f_AWID_7(h2f_AWID_7),
	.h2f_AWID_8(h2f_AWID_8),
	.h2f_AWID_9(h2f_AWID_9),
	.h2f_AWID_10(h2f_AWID_10),
	.h2f_AWID_11(h2f_AWID_11),
	.h2f_AWSIZE_0(h2f_AWSIZE_0),
	.h2f_AWSIZE_1(h2f_AWSIZE_1),
	.h2f_AWSIZE_2(h2f_AWSIZE_2),
	.h2f_WDATA_0(h2f_WDATA_0),
	.h2f_WDATA_1(h2f_WDATA_1),
	.h2f_WDATA_2(h2f_WDATA_2),
	.h2f_WDATA_3(h2f_WDATA_3),
	.h2f_WDATA_4(h2f_WDATA_4),
	.h2f_WDATA_5(h2f_WDATA_5),
	.h2f_WDATA_6(h2f_WDATA_6),
	.h2f_WDATA_7(h2f_WDATA_7),
	.h2f_WDATA_8(h2f_WDATA_8),
	.h2f_WSTRB_0(h2f_WSTRB_0),
	.h2f_WSTRB_1(h2f_WSTRB_1),
	.h2f_WSTRB_2(h2f_WSTRB_2),
	.h2f_WSTRB_3(h2f_WSTRB_3),
	.nxt_in_ready(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.nxt_in_ready1(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.saved_grant_1(\cmd_mux_005|saved_grant[1]~q ),
	.write_addr_data_both_valid(\hps_0_h2f_axi_master_agent|write_addr_data_both_valid~combout ),
	.out_data_5(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[5]~1_combout ),
	.Equal5(\router|Equal5~0_combout ),
	.Equal15(\router|Equal15~0_combout ),
	.saved_grant_0(\cmd_mux_005|saved_grant[0]~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.Equal51(\router|Equal5~1_combout ),
	.src5_valid(\cmd_demux|src5_valid~0_combout ),
	.src5_valid1(\cmd_demux|src5_valid~1_combout ),
	.cmd_src_valid_5(\hps_0_h2f_axi_master_rd_limiter|cmd_src_valid[5]~0_combout ),
	.src_valid(\cmd_mux_005|src_valid~1_combout ),
	.src_data_87(\cmd_mux_005|src_data[87]~combout ),
	.src_data_88(\cmd_mux_005|src_data[88]~combout ),
	.src_valid1(\cmd_mux_005|src_valid~2_combout ),
	.src_data_35(\cmd_mux_005|src_data[35]~combout ),
	.src_data_34(\cmd_mux_005|src_data[34]~combout ),
	.src_data_33(\cmd_mux_005|src_data[33]~combout ),
	.src_data_32(\cmd_mux_005|src_data[32]~combout ),
	.src_payload_0(\cmd_mux_005|src_payload[0]~combout ),
	.src5_valid2(\cmd_demux|src5_valid~2_combout ),
	.Selector3(\hps_0_h2f_axi_master_agent|Selector3~0_combout ),
	.Selector10(\hps_0_h2f_axi_master_agent|Selector10~1_combout ),
	.Selector4(\hps_0_h2f_axi_master_agent|Selector4~1_combout ),
	.Selector11(\hps_0_h2f_axi_master_agent|Selector11~1_combout ),
	.src_payload(\cmd_mux_005|src_payload~0_combout ),
	.src_data_82(\cmd_mux_005|src_data[82]~combout ),
	.src_data_81(\cmd_mux_005|src_data[81]~combout ),
	.src_payload1(\cmd_mux_005|src_payload~1_combout ),
	.src_payload2(\cmd_mux_005|src_payload~2_combout ),
	.src_payload3(\cmd_mux_005|src_payload~3_combout ),
	.src_payload4(\cmd_mux_005|src_payload~4_combout ),
	.src_payload5(\cmd_mux_005|src_payload~5_combout ),
	.src_payload6(\cmd_mux_005|src_payload~6_combout ),
	.src_payload7(\cmd_mux_005|src_payload~7_combout ),
	.src_payload8(\cmd_mux_005|src_payload~8_combout ),
	.src_data_105(\cmd_mux_005|src_data[105]~combout ),
	.src_data_106(\cmd_mux_005|src_data[106]~combout ),
	.src_data_107(\cmd_mux_005|src_data[107]~combout ),
	.src_data_108(\cmd_mux_005|src_data[108]~combout ),
	.src_data_109(\cmd_mux_005|src_data[109]~combout ),
	.src_data_110(\cmd_mux_005|src_data[110]~combout ),
	.src_data_111(\cmd_mux_005|src_data[111]~combout ),
	.src_data_112(\cmd_mux_005|src_data[112]~combout ),
	.src_data_113(\cmd_mux_005|src_data[113]~combout ),
	.src_data_114(\cmd_mux_005|src_data[114]~combout ),
	.src_data_115(\cmd_mux_005|src_data[115]~combout ),
	.src_data_116(\cmd_mux_005|src_data[116]~combout ),
	.src_data_86(\cmd_mux_005|src_data[86]~combout ),
	.Selector5(\hps_0_h2f_axi_master_agent|Selector5~1_combout ),
	.Selector12(\hps_0_h2f_axi_master_agent|Selector12~0_combout ),
	.src_data_80(\cmd_mux_005|src_data[80]~combout ),
	.Selector6(\hps_0_h2f_axi_master_agent|Selector6~0_combout ),
	.Selector13(\hps_0_h2f_axi_master_agent|Selector13~1_combout ),
	.src_data_79(\cmd_mux_005|src_data[79]~combout ),
	.clk_clk(clk_clk));

spw_babasu_spw_babasu_mm_interconnect_0_cmd_mux_4 cmd_mux_004(
	.h2f_ARVALID_0(h2f_ARVALID_0),
	.h2f_ARSIZE_0(h2f_ARSIZE_0),
	.h2f_ARSIZE_1(h2f_ARSIZE_1),
	.h2f_ARSIZE_2(h2f_ARSIZE_2),
	.has_pending_responses(\hps_0_h2f_axi_master_rd_limiter|has_pending_responses~q ),
	.saved_grant_1(\cmd_mux_004|saved_grant[1]~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.nxt_in_ready(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ),
	.Equal4(\router_001|Equal4~0_combout ),
	.last_channel_4(\hps_0_h2f_axi_master_rd_limiter|last_channel[4]~q ),
	.src_valid(\cmd_mux_004|src_valid~0_combout ),
	.src_payload(\cmd_mux_004|src_payload~0_combout ),
	.src_payload1(\cmd_mux_004|src_payload~1_combout ),
	.src_payload2(\cmd_mux_004|src_payload~2_combout ),
	.clk_clk(clk_clk));

spw_babasu_spw_babasu_mm_interconnect_0_cmd_mux_3 cmd_mux_003(
	.h2f_ARVALID_0(h2f_ARVALID_0),
	.h2f_ARSIZE_0(h2f_ARSIZE_0),
	.h2f_ARSIZE_1(h2f_ARSIZE_1),
	.h2f_ARSIZE_2(h2f_ARSIZE_2),
	.has_pending_responses(\hps_0_h2f_axi_master_rd_limiter|has_pending_responses~q ),
	.Equal3(\router_001|Equal3~0_combout ),
	.saved_grant_1(\cmd_mux_003|saved_grant[1]~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.nxt_in_ready(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.last_channel_3(\hps_0_h2f_axi_master_rd_limiter|last_channel[3]~q ),
	.src_valid(\cmd_mux_003|src_valid~0_combout ),
	.src_payload(\cmd_mux_003|src_payload~0_combout ),
	.src_payload1(\cmd_mux_003|src_payload~1_combout ),
	.src_payload2(\cmd_mux_003|src_payload~2_combout ),
	.clk_clk(clk_clk));

spw_babasu_spw_babasu_mm_interconnect_0_cmd_mux_2 cmd_mux_002(
	.h2f_WLAST_0(h2f_WLAST_0),
	.h2f_ARID_0(h2f_ARID_0),
	.h2f_ARID_1(h2f_ARID_1),
	.h2f_ARID_2(h2f_ARID_2),
	.h2f_ARID_3(h2f_ARID_3),
	.h2f_ARID_4(h2f_ARID_4),
	.h2f_ARID_5(h2f_ARID_5),
	.h2f_ARID_6(h2f_ARID_6),
	.h2f_ARID_7(h2f_ARID_7),
	.h2f_ARID_8(h2f_ARID_8),
	.h2f_ARID_9(h2f_ARID_9),
	.h2f_ARID_10(h2f_ARID_10),
	.h2f_ARID_11(h2f_ARID_11),
	.h2f_ARSIZE_0(h2f_ARSIZE_0),
	.h2f_ARSIZE_1(h2f_ARSIZE_1),
	.h2f_ARSIZE_2(h2f_ARSIZE_2),
	.h2f_AWID_0(h2f_AWID_0),
	.h2f_AWID_1(h2f_AWID_1),
	.h2f_AWID_2(h2f_AWID_2),
	.h2f_AWID_3(h2f_AWID_3),
	.h2f_AWID_4(h2f_AWID_4),
	.h2f_AWID_5(h2f_AWID_5),
	.h2f_AWID_6(h2f_AWID_6),
	.h2f_AWID_7(h2f_AWID_7),
	.h2f_AWID_8(h2f_AWID_8),
	.h2f_AWID_9(h2f_AWID_9),
	.h2f_AWID_10(h2f_AWID_10),
	.h2f_AWID_11(h2f_AWID_11),
	.h2f_AWSIZE_0(h2f_AWSIZE_0),
	.h2f_AWSIZE_1(h2f_AWSIZE_1),
	.h2f_AWSIZE_2(h2f_AWSIZE_2),
	.h2f_WDATA_0(h2f_WDATA_0),
	.h2f_WSTRB_0(h2f_WSTRB_0),
	.h2f_WSTRB_1(h2f_WSTRB_1),
	.h2f_WSTRB_2(h2f_WSTRB_2),
	.h2f_WSTRB_3(h2f_WSTRB_3),
	.nxt_in_ready(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.nxt_in_ready1(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.saved_grant_1(\cmd_mux_002|saved_grant[1]~q ),
	.write_addr_data_both_valid(\hps_0_h2f_axi_master_agent|write_addr_data_both_valid~combout ),
	.out_data_4(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[4]~2_combout ),
	.Equal14(\router|Equal14~0_combout ),
	.Equal16(\router|Equal16~0_combout ),
	.saved_grant_0(\cmd_mux_002|saved_grant[0]~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.Equal141(\router|Equal14~1_combout ),
	.src2_valid(\cmd_demux|src2_valid~0_combout ),
	.src2_valid1(\cmd_demux|src2_valid~1_combout ),
	.src_channel_2(\router_001|src_channel[2]~4_combout ),
	.src2_valid2(\cmd_demux_001|src2_valid~0_combout ),
	.src_valid(\cmd_mux_002|src_valid~0_combout ),
	.src_data_87(\cmd_mux_002|src_data[87]~combout ),
	.src_data_88(\cmd_mux_002|src_data[88]~combout ),
	.src_valid1(\cmd_mux_002|src_valid~1_combout ),
	.src_data_35(\cmd_mux_002|src_data[35]~combout ),
	.src_data_34(\cmd_mux_002|src_data[34]~combout ),
	.src_data_33(\cmd_mux_002|src_data[33]~combout ),
	.src_data_32(\cmd_mux_002|src_data[32]~combout ),
	.src_payload_0(\cmd_mux_002|src_payload[0]~combout ),
	.src2_valid3(\cmd_demux|src2_valid~2_combout ),
	.src2_valid4(\cmd_demux_001|src2_valid~1_combout ),
	.src_payload(\cmd_mux_002|src_payload~0_combout ),
	.Selector3(\hps_0_h2f_axi_master_agent|Selector3~0_combout ),
	.Selector10(\hps_0_h2f_axi_master_agent|Selector10~1_combout ),
	.src_data_82(\cmd_mux_002|src_data[82]~combout ),
	.Selector4(\hps_0_h2f_axi_master_agent|Selector4~1_combout ),
	.Selector11(\hps_0_h2f_axi_master_agent|Selector11~1_combout ),
	.src_data_81(\cmd_mux_002|src_data[81]~combout ),
	.src_data_105(\cmd_mux_002|src_data[105]~combout ),
	.src_data_106(\cmd_mux_002|src_data[106]~combout ),
	.src_data_107(\cmd_mux_002|src_data[107]~combout ),
	.src_data_108(\cmd_mux_002|src_data[108]~combout ),
	.src_data_109(\cmd_mux_002|src_data[109]~combout ),
	.src_data_110(\cmd_mux_002|src_data[110]~combout ),
	.src_data_111(\cmd_mux_002|src_data[111]~combout ),
	.src_data_112(\cmd_mux_002|src_data[112]~combout ),
	.src_data_113(\cmd_mux_002|src_data[113]~combout ),
	.src_data_114(\cmd_mux_002|src_data[114]~combout ),
	.src_data_115(\cmd_mux_002|src_data[115]~combout ),
	.src_data_116(\cmd_mux_002|src_data[116]~combout ),
	.src_data_86(\cmd_mux_002|src_data[86]~combout ),
	.Selector5(\hps_0_h2f_axi_master_agent|Selector5~1_combout ),
	.Selector12(\hps_0_h2f_axi_master_agent|Selector12~0_combout ),
	.src_data_80(\cmd_mux_002|src_data[80]~combout ),
	.Selector6(\hps_0_h2f_axi_master_agent|Selector6~0_combout ),
	.Selector13(\hps_0_h2f_axi_master_agent|Selector13~1_combout ),
	.src_data_79(\cmd_mux_002|src_data[79]~combout ),
	.clk_clk(clk_clk));

spw_babasu_spw_babasu_mm_interconnect_0_cmd_mux_1 cmd_mux_001(
	.h2f_ARVALID_0(h2f_ARVALID_0),
	.h2f_WLAST_0(h2f_WLAST_0),
	.h2f_ARID_0(h2f_ARID_0),
	.h2f_ARID_1(h2f_ARID_1),
	.h2f_ARID_2(h2f_ARID_2),
	.h2f_ARID_3(h2f_ARID_3),
	.h2f_ARID_4(h2f_ARID_4),
	.h2f_ARID_5(h2f_ARID_5),
	.h2f_ARID_6(h2f_ARID_6),
	.h2f_ARID_7(h2f_ARID_7),
	.h2f_ARID_8(h2f_ARID_8),
	.h2f_ARID_9(h2f_ARID_9),
	.h2f_ARID_10(h2f_ARID_10),
	.h2f_ARID_11(h2f_ARID_11),
	.h2f_ARSIZE_0(h2f_ARSIZE_0),
	.h2f_ARSIZE_1(h2f_ARSIZE_1),
	.h2f_ARSIZE_2(h2f_ARSIZE_2),
	.h2f_AWID_0(h2f_AWID_0),
	.h2f_AWID_1(h2f_AWID_1),
	.h2f_AWID_2(h2f_AWID_2),
	.h2f_AWID_3(h2f_AWID_3),
	.h2f_AWID_4(h2f_AWID_4),
	.h2f_AWID_5(h2f_AWID_5),
	.h2f_AWID_6(h2f_AWID_6),
	.h2f_AWID_7(h2f_AWID_7),
	.h2f_AWID_8(h2f_AWID_8),
	.h2f_AWID_9(h2f_AWID_9),
	.h2f_AWID_10(h2f_AWID_10),
	.h2f_AWID_11(h2f_AWID_11),
	.h2f_AWSIZE_0(h2f_AWSIZE_0),
	.h2f_AWSIZE_1(h2f_AWSIZE_1),
	.h2f_AWSIZE_2(h2f_AWSIZE_2),
	.h2f_WDATA_0(h2f_WDATA_0),
	.h2f_WSTRB_0(h2f_WSTRB_0),
	.h2f_WSTRB_1(h2f_WSTRB_1),
	.h2f_WSTRB_2(h2f_WSTRB_2),
	.h2f_WSTRB_3(h2f_WSTRB_3),
	.nxt_in_ready(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.has_pending_responses(\hps_0_h2f_axi_master_rd_limiter|has_pending_responses~q ),
	.nxt_in_ready1(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.saved_grant_1(\cmd_mux_001|saved_grant[1]~q ),
	.src_channel_1(\router_001|src_channel[1]~1_combout ),
	.write_addr_data_both_valid(\hps_0_h2f_axi_master_agent|write_addr_data_both_valid~combout ),
	.out_data_5(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[5]~1_combout ),
	.Equal16(\router|Equal16~0_combout ),
	.Equal15(\router|Equal15~0_combout ),
	.saved_grant_0(\cmd_mux_001|saved_grant[0]~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.Equal5(\router|Equal5~1_combout ),
	.src1_valid(\cmd_demux|src1_valid~0_combout ),
	.src1_valid1(\cmd_demux|src1_valid~1_combout ),
	.last_channel_1(\hps_0_h2f_axi_master_rd_limiter|last_channel[1]~q ),
	.src_valid(\cmd_mux_001|src_valid~0_combout ),
	.src_data_87(\cmd_mux_001|src_data[87]~combout ),
	.src_data_88(\cmd_mux_001|src_data[88]~combout ),
	.src_valid1(\cmd_mux_001|src_valid~1_combout ),
	.src_data_35(\cmd_mux_001|src_data[35]~combout ),
	.src_data_34(\cmd_mux_001|src_data[34]~combout ),
	.src_data_33(\cmd_mux_001|src_data[33]~combout ),
	.src_data_32(\cmd_mux_001|src_data[32]~combout ),
	.src_payload_0(\cmd_mux_001|src_payload[0]~combout ),
	.src1_valid2(\cmd_demux|src1_valid~2_combout ),
	.src1_valid3(\cmd_demux_001|src1_valid~0_combout ),
	.Selector3(\hps_0_h2f_axi_master_agent|Selector3~0_combout ),
	.Selector10(\hps_0_h2f_axi_master_agent|Selector10~1_combout ),
	.Selector4(\hps_0_h2f_axi_master_agent|Selector4~1_combout ),
	.Selector11(\hps_0_h2f_axi_master_agent|Selector11~1_combout ),
	.src_payload(\cmd_mux_001|src_payload~0_combout ),
	.src_data_82(\cmd_mux_001|src_data[82]~combout ),
	.src_data_81(\cmd_mux_001|src_data[81]~combout ),
	.src_data_105(\cmd_mux_001|src_data[105]~combout ),
	.src_data_106(\cmd_mux_001|src_data[106]~combout ),
	.src_data_107(\cmd_mux_001|src_data[107]~combout ),
	.src_data_108(\cmd_mux_001|src_data[108]~combout ),
	.src_data_109(\cmd_mux_001|src_data[109]~combout ),
	.src_data_110(\cmd_mux_001|src_data[110]~combout ),
	.src_data_111(\cmd_mux_001|src_data[111]~combout ),
	.src_data_112(\cmd_mux_001|src_data[112]~combout ),
	.src_data_113(\cmd_mux_001|src_data[113]~combout ),
	.src_data_114(\cmd_mux_001|src_data[114]~combout ),
	.src_data_115(\cmd_mux_001|src_data[115]~combout ),
	.src_data_116(\cmd_mux_001|src_data[116]~combout ),
	.src_data_86(\cmd_mux_001|src_data[86]~combout ),
	.Selector5(\hps_0_h2f_axi_master_agent|Selector5~1_combout ),
	.Selector12(\hps_0_h2f_axi_master_agent|Selector12~0_combout ),
	.src_data_80(\cmd_mux_001|src_data[80]~combout ),
	.Selector6(\hps_0_h2f_axi_master_agent|Selector6~0_combout ),
	.Selector13(\hps_0_h2f_axi_master_agent|Selector13~1_combout ),
	.src_data_79(\cmd_mux_001|src_data[79]~combout ),
	.clk_clk(clk_clk));

spw_babasu_spw_babasu_mm_interconnect_0_rsp_demux_5 rsp_demux_005(
	.h2f_BREADY_0(h2f_BREADY_0),
	.h2f_RREADY_0(h2f_RREADY_0),
	.read_latency_shift_reg_0(\data_i_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\data_i_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_129_0(\data_i_s1_agent_rsp_fifo|mem[0][129]~q ),
	.mem_used_01(\data_i_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_68_0(\data_i_s1_agent_rsp_fifo|mem[0][68]~q ),
	.mem_66_0(\data_i_s1_agent_rsp_fifo|mem[0][66]~q ),
	.src0_valid1(\rsp_demux_005|src0_valid~combout ),
	.src1_valid(\rsp_demux_005|src1_valid~0_combout ),
	.WideOr0(\rsp_demux_005|WideOr0~0_combout ));

spw_babasu_spw_babasu_mm_interconnect_0_rsp_demux_2 rsp_demux_002(
	.h2f_BREADY_0(h2f_BREADY_0),
	.h2f_RREADY_0(h2f_RREADY_0),
	.read_latency_shift_reg_0(\autostart_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\autostart_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_129_0(\autostart_s1_agent_rsp_fifo|mem[0][129]~q ),
	.mem_used_01(\autostart_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_68_0(\autostart_s1_agent_rsp_fifo|mem[0][68]~q ),
	.mem_66_0(\autostart_s1_agent_rsp_fifo|mem[0][66]~q ),
	.src0_valid1(\rsp_demux_002|src0_valid~combout ),
	.src1_valid(\rsp_demux_002|src1_valid~0_combout ),
	.WideOr0(\rsp_demux_002|WideOr0~0_combout ));

spw_babasu_spw_babasu_mm_interconnect_0_rsp_demux_1 rsp_demux_001(
	.h2f_BREADY_0(h2f_BREADY_0),
	.h2f_RREADY_0(h2f_RREADY_0),
	.read_latency_shift_reg_0(\link_disable_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\link_disable_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_129_0(\link_disable_s1_agent_rsp_fifo|mem[0][129]~q ),
	.mem_used_01(\link_disable_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_68_0(\link_disable_s1_agent_rsp_fifo|mem[0][68]~q ),
	.mem_66_0(\link_disable_s1_agent_rsp_fifo|mem[0][66]~q ),
	.src0_valid1(\rsp_demux_001|src0_valid~combout ),
	.src1_valid(\rsp_demux_001|src1_valid~0_combout ),
	.WideOr0(\rsp_demux_001|WideOr0~0_combout ));

spw_babasu_spw_babasu_mm_interconnect_0_rsp_demux rsp_demux(
	.h2f_BREADY_0(h2f_BREADY_0),
	.h2f_RREADY_0(h2f_RREADY_0),
	.read_latency_shift_reg_0(\link_start_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\link_start_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_129_0(\link_start_s1_agent_rsp_fifo|mem[0][129]~q ),
	.mem_used_01(\link_start_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_68_0(\link_start_s1_agent_rsp_fifo|mem[0][68]~q ),
	.mem_66_0(\link_start_s1_agent_rsp_fifo|mem[0][66]~q ),
	.src0_valid1(\rsp_demux|src0_valid~combout ),
	.src1_valid(\rsp_demux|src1_valid~0_combout ),
	.WideOr0(\rsp_demux|WideOr0~0_combout ));

spw_babasu_spw_babasu_mm_interconnect_0_cmd_mux_16 cmd_mux_016(
	.h2f_WLAST_0(h2f_WLAST_0),
	.h2f_ARID_0(h2f_ARID_0),
	.h2f_ARID_1(h2f_ARID_1),
	.h2f_ARID_2(h2f_ARID_2),
	.h2f_ARID_3(h2f_ARID_3),
	.h2f_ARID_4(h2f_ARID_4),
	.h2f_ARID_5(h2f_ARID_5),
	.h2f_ARID_6(h2f_ARID_6),
	.h2f_ARID_7(h2f_ARID_7),
	.h2f_ARID_8(h2f_ARID_8),
	.h2f_ARID_9(h2f_ARID_9),
	.h2f_ARID_10(h2f_ARID_10),
	.h2f_ARID_11(h2f_ARID_11),
	.h2f_ARSIZE_0(h2f_ARSIZE_0),
	.h2f_ARSIZE_1(h2f_ARSIZE_1),
	.h2f_ARSIZE_2(h2f_ARSIZE_2),
	.h2f_AWID_0(h2f_AWID_0),
	.h2f_AWID_1(h2f_AWID_1),
	.h2f_AWID_2(h2f_AWID_2),
	.h2f_AWID_3(h2f_AWID_3),
	.h2f_AWID_4(h2f_AWID_4),
	.h2f_AWID_5(h2f_AWID_5),
	.h2f_AWID_6(h2f_AWID_6),
	.h2f_AWID_7(h2f_AWID_7),
	.h2f_AWID_8(h2f_AWID_8),
	.h2f_AWID_9(h2f_AWID_9),
	.h2f_AWID_10(h2f_AWID_10),
	.h2f_AWID_11(h2f_AWID_11),
	.h2f_AWSIZE_0(h2f_AWSIZE_0),
	.h2f_AWSIZE_1(h2f_AWSIZE_1),
	.h2f_AWSIZE_2(h2f_AWSIZE_2),
	.h2f_WDATA_0(h2f_WDATA_0),
	.h2f_WSTRB_0(h2f_WSTRB_0),
	.h2f_WSTRB_1(h2f_WSTRB_1),
	.h2f_WSTRB_2(h2f_WSTRB_2),
	.h2f_WSTRB_3(h2f_WSTRB_3),
	.nxt_in_ready(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ),
	.nxt_in_ready1(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.Equal16(\router_001|Equal16~0_combout ),
	.saved_grant_1(\cmd_mux_016|saved_grant[1]~q ),
	.write_addr_data_both_valid(\hps_0_h2f_axi_master_agent|write_addr_data_both_valid~combout ),
	.out_data_4(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[4]~2_combout ),
	.Equal161(\router|Equal16~0_combout ),
	.Equal162(\router|Equal16~1_combout ),
	.saved_grant_0(\cmd_mux_016|saved_grant[0]~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.src16_valid(\cmd_demux|src16_valid~0_combout ),
	.src16_valid1(\cmd_demux|src16_valid~1_combout ),
	.src16_valid2(\cmd_demux_001|src16_valid~0_combout ),
	.src_valid(\cmd_mux_016|src_valid~0_combout ),
	.src_valid1(\cmd_mux_016|src_valid~1_combout ),
	.src16_valid3(\cmd_demux|src16_valid~2_combout ),
	.WideOr11(\cmd_mux_016|WideOr1~combout ),
	.src_data_87(\cmd_mux_016|src_data[87]~combout ),
	.src_data_88(\cmd_mux_016|src_data[88]~combout ),
	.src_data_35(\cmd_mux_016|src_data[35]~combout ),
	.src_data_34(\cmd_mux_016|src_data[34]~combout ),
	.src_data_33(\cmd_mux_016|src_data[33]~combout ),
	.src_data_32(\cmd_mux_016|src_data[32]~combout ),
	.src_payload_0(\cmd_mux_016|src_payload[0]~combout ),
	.src16_valid4(\cmd_demux_001|src16_valid~1_combout ),
	.Selector3(\hps_0_h2f_axi_master_agent|Selector3~0_combout ),
	.Selector10(\hps_0_h2f_axi_master_agent|Selector10~1_combout ),
	.Selector4(\hps_0_h2f_axi_master_agent|Selector4~1_combout ),
	.Selector11(\hps_0_h2f_axi_master_agent|Selector11~1_combout ),
	.src_payload(\cmd_mux_016|src_payload~0_combout ),
	.src_data_82(\cmd_mux_016|src_data[82]~combout ),
	.src_data_81(\cmd_mux_016|src_data[81]~combout ),
	.src_data_105(\cmd_mux_016|src_data[105]~combout ),
	.src_data_106(\cmd_mux_016|src_data[106]~combout ),
	.src_data_107(\cmd_mux_016|src_data[107]~combout ),
	.src_data_108(\cmd_mux_016|src_data[108]~combout ),
	.src_data_109(\cmd_mux_016|src_data[109]~combout ),
	.src_data_110(\cmd_mux_016|src_data[110]~combout ),
	.src_data_111(\cmd_mux_016|src_data[111]~combout ),
	.src_data_112(\cmd_mux_016|src_data[112]~combout ),
	.src_data_113(\cmd_mux_016|src_data[113]~combout ),
	.src_data_114(\cmd_mux_016|src_data[114]~combout ),
	.src_data_115(\cmd_mux_016|src_data[115]~combout ),
	.src_data_116(\cmd_mux_016|src_data[116]~combout ),
	.src_data_86(\cmd_mux_016|src_data[86]~combout ),
	.Selector5(\hps_0_h2f_axi_master_agent|Selector5~1_combout ),
	.Selector12(\hps_0_h2f_axi_master_agent|Selector12~0_combout ),
	.src_data_80(\cmd_mux_016|src_data[80]~combout ),
	.Selector6(\hps_0_h2f_axi_master_agent|Selector6~0_combout ),
	.Selector13(\hps_0_h2f_axi_master_agent|Selector13~1_combout ),
	.src_data_79(\cmd_mux_016|src_data[79]~combout ),
	.clk_clk(clk_clk));

spw_babasu_spw_babasu_mm_interconnect_0_cmd_mux_15 cmd_mux_015(
	.h2f_WLAST_0(h2f_WLAST_0),
	.h2f_ARID_0(h2f_ARID_0),
	.h2f_ARID_1(h2f_ARID_1),
	.h2f_ARID_2(h2f_ARID_2),
	.h2f_ARID_3(h2f_ARID_3),
	.h2f_ARID_4(h2f_ARID_4),
	.h2f_ARID_5(h2f_ARID_5),
	.h2f_ARID_6(h2f_ARID_6),
	.h2f_ARID_7(h2f_ARID_7),
	.h2f_ARID_8(h2f_ARID_8),
	.h2f_ARID_9(h2f_ARID_9),
	.h2f_ARID_10(h2f_ARID_10),
	.h2f_ARID_11(h2f_ARID_11),
	.h2f_ARSIZE_0(h2f_ARSIZE_0),
	.h2f_ARSIZE_1(h2f_ARSIZE_1),
	.h2f_ARSIZE_2(h2f_ARSIZE_2),
	.h2f_AWID_0(h2f_AWID_0),
	.h2f_AWID_1(h2f_AWID_1),
	.h2f_AWID_2(h2f_AWID_2),
	.h2f_AWID_3(h2f_AWID_3),
	.h2f_AWID_4(h2f_AWID_4),
	.h2f_AWID_5(h2f_AWID_5),
	.h2f_AWID_6(h2f_AWID_6),
	.h2f_AWID_7(h2f_AWID_7),
	.h2f_AWID_8(h2f_AWID_8),
	.h2f_AWID_9(h2f_AWID_9),
	.h2f_AWID_10(h2f_AWID_10),
	.h2f_AWID_11(h2f_AWID_11),
	.h2f_AWSIZE_0(h2f_AWSIZE_0),
	.h2f_AWSIZE_1(h2f_AWSIZE_1),
	.h2f_AWSIZE_2(h2f_AWSIZE_2),
	.h2f_WDATA_0(h2f_WDATA_0),
	.h2f_WDATA_1(h2f_WDATA_1),
	.h2f_WDATA_2(h2f_WDATA_2),
	.h2f_WDATA_3(h2f_WDATA_3),
	.h2f_WDATA_4(h2f_WDATA_4),
	.h2f_WDATA_5(h2f_WDATA_5),
	.h2f_WDATA_6(h2f_WDATA_6),
	.h2f_WSTRB_0(h2f_WSTRB_0),
	.h2f_WSTRB_1(h2f_WSTRB_1),
	.h2f_WSTRB_2(h2f_WSTRB_2),
	.h2f_WSTRB_3(h2f_WSTRB_3),
	.nxt_in_ready(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.nxt_in_ready1(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.saved_grant_1(\cmd_mux_015|saved_grant[1]~q ),
	.Equal15(\router_001|Equal15~0_combout ),
	.write_addr_data_both_valid(\hps_0_h2f_axi_master_agent|write_addr_data_both_valid~combout ),
	.out_data_5(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[5]~1_combout ),
	.Equal13(\router|Equal13~0_combout ),
	.Equal151(\router|Equal15~0_combout ),
	.saved_grant_0(\cmd_mux_015|saved_grant[0]~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.Equal152(\router|Equal15~1_combout ),
	.src15_valid(\cmd_demux|src15_valid~0_combout ),
	.src15_valid1(\cmd_demux|src15_valid~1_combout ),
	.src15_valid2(\cmd_demux_001|src15_valid~0_combout ),
	.src_valid(\cmd_mux_015|src_valid~0_combout ),
	.src_data_87(\cmd_mux_015|src_data[87]~combout ),
	.src_data_88(\cmd_mux_015|src_data[88]~combout ),
	.src_valid1(\cmd_mux_015|src_valid~1_combout ),
	.src_data_35(\cmd_mux_015|src_data[35]~combout ),
	.src_data_34(\cmd_mux_015|src_data[34]~combout ),
	.src_data_33(\cmd_mux_015|src_data[33]~combout ),
	.src_data_32(\cmd_mux_015|src_data[32]~combout ),
	.src_payload_0(\cmd_mux_015|src_payload[0]~combout ),
	.src15_valid3(\cmd_demux|src15_valid~2_combout ),
	.src15_valid4(\cmd_demux_001|src15_valid~1_combout ),
	.Selector3(\hps_0_h2f_axi_master_agent|Selector3~0_combout ),
	.Selector10(\hps_0_h2f_axi_master_agent|Selector10~1_combout ),
	.Selector4(\hps_0_h2f_axi_master_agent|Selector4~1_combout ),
	.Selector11(\hps_0_h2f_axi_master_agent|Selector11~1_combout ),
	.src_payload(\cmd_mux_015|src_payload~0_combout ),
	.src_data_82(\cmd_mux_015|src_data[82]~combout ),
	.src_data_81(\cmd_mux_015|src_data[81]~combout ),
	.src_payload1(\cmd_mux_015|src_payload~1_combout ),
	.src_payload2(\cmd_mux_015|src_payload~2_combout ),
	.src_payload3(\cmd_mux_015|src_payload~3_combout ),
	.src_payload4(\cmd_mux_015|src_payload~4_combout ),
	.src_payload5(\cmd_mux_015|src_payload~5_combout ),
	.src_payload6(\cmd_mux_015|src_payload~6_combout ),
	.src_data_105(\cmd_mux_015|src_data[105]~combout ),
	.src_data_106(\cmd_mux_015|src_data[106]~combout ),
	.src_data_107(\cmd_mux_015|src_data[107]~combout ),
	.src_data_108(\cmd_mux_015|src_data[108]~combout ),
	.src_data_109(\cmd_mux_015|src_data[109]~combout ),
	.src_data_110(\cmd_mux_015|src_data[110]~combout ),
	.src_data_111(\cmd_mux_015|src_data[111]~combout ),
	.src_data_112(\cmd_mux_015|src_data[112]~combout ),
	.src_data_113(\cmd_mux_015|src_data[113]~combout ),
	.src_data_114(\cmd_mux_015|src_data[114]~combout ),
	.src_data_115(\cmd_mux_015|src_data[115]~combout ),
	.src_data_116(\cmd_mux_015|src_data[116]~combout ),
	.src_data_86(\cmd_mux_015|src_data[86]~combout ),
	.Selector5(\hps_0_h2f_axi_master_agent|Selector5~1_combout ),
	.Selector12(\hps_0_h2f_axi_master_agent|Selector12~0_combout ),
	.src_data_80(\cmd_mux_015|src_data[80]~combout ),
	.Selector6(\hps_0_h2f_axi_master_agent|Selector6~0_combout ),
	.Selector13(\hps_0_h2f_axi_master_agent|Selector13~1_combout ),
	.src_data_79(\cmd_mux_015|src_data[79]~combout ),
	.clk_clk(clk_clk));

spw_babasu_spw_babasu_mm_interconnect_0_cmd_mux_14 cmd_mux_014(
	.h2f_WLAST_0(h2f_WLAST_0),
	.h2f_ARID_0(h2f_ARID_0),
	.h2f_ARID_1(h2f_ARID_1),
	.h2f_ARID_2(h2f_ARID_2),
	.h2f_ARID_3(h2f_ARID_3),
	.h2f_ARID_4(h2f_ARID_4),
	.h2f_ARID_5(h2f_ARID_5),
	.h2f_ARID_6(h2f_ARID_6),
	.h2f_ARID_7(h2f_ARID_7),
	.h2f_ARID_8(h2f_ARID_8),
	.h2f_ARID_9(h2f_ARID_9),
	.h2f_ARID_10(h2f_ARID_10),
	.h2f_ARID_11(h2f_ARID_11),
	.h2f_ARSIZE_0(h2f_ARSIZE_0),
	.h2f_ARSIZE_1(h2f_ARSIZE_1),
	.h2f_ARSIZE_2(h2f_ARSIZE_2),
	.h2f_AWID_0(h2f_AWID_0),
	.h2f_AWID_1(h2f_AWID_1),
	.h2f_AWID_2(h2f_AWID_2),
	.h2f_AWID_3(h2f_AWID_3),
	.h2f_AWID_4(h2f_AWID_4),
	.h2f_AWID_5(h2f_AWID_5),
	.h2f_AWID_6(h2f_AWID_6),
	.h2f_AWID_7(h2f_AWID_7),
	.h2f_AWID_8(h2f_AWID_8),
	.h2f_AWID_9(h2f_AWID_9),
	.h2f_AWID_10(h2f_AWID_10),
	.h2f_AWID_11(h2f_AWID_11),
	.h2f_AWSIZE_0(h2f_AWSIZE_0),
	.h2f_AWSIZE_1(h2f_AWSIZE_1),
	.h2f_AWSIZE_2(h2f_AWSIZE_2),
	.h2f_WDATA_0(h2f_WDATA_0),
	.h2f_WDATA_1(h2f_WDATA_1),
	.h2f_WDATA_2(h2f_WDATA_2),
	.h2f_WDATA_3(h2f_WDATA_3),
	.h2f_WDATA_4(h2f_WDATA_4),
	.h2f_WDATA_5(h2f_WDATA_5),
	.h2f_WDATA_6(h2f_WDATA_6),
	.h2f_WDATA_7(h2f_WDATA_7),
	.h2f_WSTRB_0(h2f_WSTRB_0),
	.h2f_WSTRB_1(h2f_WSTRB_1),
	.h2f_WSTRB_2(h2f_WSTRB_2),
	.h2f_WSTRB_3(h2f_WSTRB_3),
	.nxt_in_ready(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.nxt_in_ready1(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.saved_grant_1(\cmd_mux_014|saved_grant[1]~q ),
	.Equal14(\router_001|Equal14~0_combout ),
	.write_addr_data_both_valid(\hps_0_h2f_axi_master_agent|write_addr_data_both_valid~combout ),
	.out_data_4(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[4]~2_combout ),
	.Equal141(\router|Equal14~0_combout ),
	.Equal13(\router|Equal13~0_combout ),
	.saved_grant_0(\cmd_mux_014|saved_grant[0]~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.Equal142(\router|Equal14~1_combout ),
	.src14_valid(\cmd_demux|src14_valid~0_combout ),
	.src14_valid1(\cmd_demux|src14_valid~1_combout ),
	.src14_valid2(\cmd_demux_001|src14_valid~0_combout ),
	.src_valid(\cmd_mux_014|src_valid~0_combout ),
	.src_data_87(\cmd_mux_014|src_data[87]~combout ),
	.src_data_88(\cmd_mux_014|src_data[88]~combout ),
	.src_valid1(\cmd_mux_014|src_valid~1_combout ),
	.src_data_35(\cmd_mux_014|src_data[35]~combout ),
	.src_data_34(\cmd_mux_014|src_data[34]~combout ),
	.src_data_33(\cmd_mux_014|src_data[33]~combout ),
	.src_data_32(\cmd_mux_014|src_data[32]~combout ),
	.src_payload_0(\cmd_mux_014|src_payload[0]~combout ),
	.src14_valid3(\cmd_demux|src14_valid~2_combout ),
	.src14_valid4(\cmd_demux_001|src14_valid~1_combout ),
	.Selector3(\hps_0_h2f_axi_master_agent|Selector3~0_combout ),
	.Selector10(\hps_0_h2f_axi_master_agent|Selector10~1_combout ),
	.Selector4(\hps_0_h2f_axi_master_agent|Selector4~1_combout ),
	.Selector11(\hps_0_h2f_axi_master_agent|Selector11~1_combout ),
	.src_payload(\cmd_mux_014|src_payload~0_combout ),
	.src_data_82(\cmd_mux_014|src_data[82]~combout ),
	.src_data_81(\cmd_mux_014|src_data[81]~combout ),
	.src_payload1(\cmd_mux_014|src_payload~1_combout ),
	.src_payload2(\cmd_mux_014|src_payload~2_combout ),
	.src_payload3(\cmd_mux_014|src_payload~3_combout ),
	.src_payload4(\cmd_mux_014|src_payload~4_combout ),
	.src_payload5(\cmd_mux_014|src_payload~5_combout ),
	.src_payload6(\cmd_mux_014|src_payload~6_combout ),
	.src_payload7(\cmd_mux_014|src_payload~7_combout ),
	.src_data_105(\cmd_mux_014|src_data[105]~combout ),
	.src_data_106(\cmd_mux_014|src_data[106]~combout ),
	.src_data_107(\cmd_mux_014|src_data[107]~combout ),
	.src_data_108(\cmd_mux_014|src_data[108]~combout ),
	.src_data_109(\cmd_mux_014|src_data[109]~combout ),
	.src_data_110(\cmd_mux_014|src_data[110]~combout ),
	.src_data_111(\cmd_mux_014|src_data[111]~combout ),
	.src_data_112(\cmd_mux_014|src_data[112]~combout ),
	.src_data_113(\cmd_mux_014|src_data[113]~combout ),
	.src_data_114(\cmd_mux_014|src_data[114]~combout ),
	.src_data_115(\cmd_mux_014|src_data[115]~combout ),
	.src_data_116(\cmd_mux_014|src_data[116]~combout ),
	.src_data_86(\cmd_mux_014|src_data[86]~combout ),
	.Selector5(\hps_0_h2f_axi_master_agent|Selector5~1_combout ),
	.Selector12(\hps_0_h2f_axi_master_agent|Selector12~0_combout ),
	.src_data_80(\cmd_mux_014|src_data[80]~combout ),
	.Selector6(\hps_0_h2f_axi_master_agent|Selector6~0_combout ),
	.Selector13(\hps_0_h2f_axi_master_agent|Selector13~1_combout ),
	.src_data_79(\cmd_mux_014|src_data[79]~combout ),
	.clk_clk(clk_clk));

spw_babasu_spw_babasu_mm_interconnect_0_cmd_mux_13 cmd_mux_013(
	.h2f_ARVALID_0(h2f_ARVALID_0),
	.h2f_WLAST_0(h2f_WLAST_0),
	.h2f_ARADDR_4(h2f_ARADDR_4),
	.h2f_ARADDR_5(h2f_ARADDR_5),
	.h2f_ARADDR_6(h2f_ARADDR_6),
	.h2f_ARADDR_7(h2f_ARADDR_7),
	.h2f_ARADDR_8(h2f_ARADDR_8),
	.h2f_ARID_0(h2f_ARID_0),
	.h2f_ARID_1(h2f_ARID_1),
	.h2f_ARID_2(h2f_ARID_2),
	.h2f_ARID_3(h2f_ARID_3),
	.h2f_ARID_4(h2f_ARID_4),
	.h2f_ARID_5(h2f_ARID_5),
	.h2f_ARID_6(h2f_ARID_6),
	.h2f_ARID_7(h2f_ARID_7),
	.h2f_ARID_8(h2f_ARID_8),
	.h2f_ARID_9(h2f_ARID_9),
	.h2f_ARID_10(h2f_ARID_10),
	.h2f_ARID_11(h2f_ARID_11),
	.h2f_ARSIZE_0(h2f_ARSIZE_0),
	.h2f_ARSIZE_1(h2f_ARSIZE_1),
	.h2f_ARSIZE_2(h2f_ARSIZE_2),
	.h2f_AWID_0(h2f_AWID_0),
	.h2f_AWID_1(h2f_AWID_1),
	.h2f_AWID_2(h2f_AWID_2),
	.h2f_AWID_3(h2f_AWID_3),
	.h2f_AWID_4(h2f_AWID_4),
	.h2f_AWID_5(h2f_AWID_5),
	.h2f_AWID_6(h2f_AWID_6),
	.h2f_AWID_7(h2f_AWID_7),
	.h2f_AWID_8(h2f_AWID_8),
	.h2f_AWID_9(h2f_AWID_9),
	.h2f_AWID_10(h2f_AWID_10),
	.h2f_AWID_11(h2f_AWID_11),
	.h2f_AWSIZE_0(h2f_AWSIZE_0),
	.h2f_AWSIZE_1(h2f_AWSIZE_1),
	.h2f_AWSIZE_2(h2f_AWSIZE_2),
	.h2f_WDATA_0(h2f_WDATA_0),
	.h2f_WSTRB_0(h2f_WSTRB_0),
	.h2f_WSTRB_1(h2f_WSTRB_1),
	.h2f_WSTRB_2(h2f_WSTRB_2),
	.h2f_WSTRB_3(h2f_WSTRB_3),
	.nxt_in_ready(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.has_pending_responses(\hps_0_h2f_axi_master_rd_limiter|has_pending_responses~q ),
	.nxt_in_ready1(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.saved_grant_1(\cmd_mux_013|saved_grant[1]~q ),
	.write_addr_data_both_valid(\hps_0_h2f_axi_master_agent|write_addr_data_both_valid~combout ),
	.out_data_5(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[5]~1_combout ),
	.Equal13(\router|Equal13~0_combout ),
	.Equal15(\router|Equal15~0_combout ),
	.saved_grant_0(\cmd_mux_013|saved_grant[0]~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.Equal5(\router|Equal5~1_combout ),
	.src13_valid(\cmd_demux|src13_valid~0_combout ),
	.src13_valid1(\cmd_demux|src13_valid~1_combout ),
	.last_channel_13(\hps_0_h2f_axi_master_rd_limiter|last_channel[13]~q ),
	.src_valid(\cmd_mux_013|src_valid~2_combout ),
	.src_data_87(\cmd_mux_013|src_data[87]~combout ),
	.src_data_88(\cmd_mux_013|src_data[88]~combout ),
	.src_valid1(\cmd_mux_013|src_valid~3_combout ),
	.src_data_35(\cmd_mux_013|src_data[35]~combout ),
	.src_data_34(\cmd_mux_013|src_data[34]~combout ),
	.src_data_33(\cmd_mux_013|src_data[33]~combout ),
	.src_data_32(\cmd_mux_013|src_data[32]~combout ),
	.src_payload_0(\cmd_mux_013|src_payload[0]~combout ),
	.src13_valid2(\cmd_demux|src13_valid~2_combout ),
	.Selector3(\hps_0_h2f_axi_master_agent|Selector3~0_combout ),
	.Selector10(\hps_0_h2f_axi_master_agent|Selector10~1_combout ),
	.Selector4(\hps_0_h2f_axi_master_agent|Selector4~1_combout ),
	.Selector11(\hps_0_h2f_axi_master_agent|Selector11~1_combout ),
	.src_payload(\cmd_mux_013|src_payload~0_combout ),
	.src_data_82(\cmd_mux_013|src_data[82]~combout ),
	.src_data_81(\cmd_mux_013|src_data[81]~combout ),
	.src_data_105(\cmd_mux_013|src_data[105]~combout ),
	.src_data_106(\cmd_mux_013|src_data[106]~combout ),
	.src_data_107(\cmd_mux_013|src_data[107]~combout ),
	.src_data_108(\cmd_mux_013|src_data[108]~combout ),
	.src_data_109(\cmd_mux_013|src_data[109]~combout ),
	.src_data_110(\cmd_mux_013|src_data[110]~combout ),
	.src_data_111(\cmd_mux_013|src_data[111]~combout ),
	.src_data_112(\cmd_mux_013|src_data[112]~combout ),
	.src_data_113(\cmd_mux_013|src_data[113]~combout ),
	.src_data_114(\cmd_mux_013|src_data[114]~combout ),
	.src_data_115(\cmd_mux_013|src_data[115]~combout ),
	.src_data_116(\cmd_mux_013|src_data[116]~combout ),
	.src_data_86(\cmd_mux_013|src_data[86]~combout ),
	.Selector5(\hps_0_h2f_axi_master_agent|Selector5~1_combout ),
	.Selector12(\hps_0_h2f_axi_master_agent|Selector12~0_combout ),
	.src_data_80(\cmd_mux_013|src_data[80]~combout ),
	.Selector6(\hps_0_h2f_axi_master_agent|Selector6~0_combout ),
	.Selector13(\hps_0_h2f_axi_master_agent|Selector13~1_combout ),
	.src_data_79(\cmd_mux_013|src_data[79]~combout ),
	.clk_clk(clk_clk));

spw_babasu_spw_babasu_mm_interconnect_0_cmd_mux_12 cmd_mux_012(
	.h2f_ARVALID_0(h2f_ARVALID_0),
	.h2f_ARADDR_4(h2f_ARADDR_4),
	.h2f_ARADDR_5(h2f_ARADDR_5),
	.h2f_ARADDR_6(h2f_ARADDR_6),
	.h2f_ARADDR_7(h2f_ARADDR_7),
	.h2f_ARADDR_8(h2f_ARADDR_8),
	.h2f_ARSIZE_0(h2f_ARSIZE_0),
	.h2f_ARSIZE_1(h2f_ARSIZE_1),
	.h2f_ARSIZE_2(h2f_ARSIZE_2),
	.has_pending_responses(\hps_0_h2f_axi_master_rd_limiter|has_pending_responses~q ),
	.saved_grant_1(\cmd_mux_012|saved_grant[1]~q ),
	.last_cycle(\cmd_mux_012|last_cycle~0_combout ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.nxt_in_ready(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.last_channel_12(\hps_0_h2f_axi_master_rd_limiter|last_channel[12]~q ),
	.src_valid(\cmd_mux_012|src_valid~0_combout ),
	.src_payload(\cmd_mux_012|src_payload~0_combout ),
	.src_payload1(\cmd_mux_012|src_payload~1_combout ),
	.src_payload2(\cmd_mux_012|src_payload~2_combout ),
	.clk_clk(clk_clk));

spw_babasu_spw_babasu_mm_interconnect_0_cmd_mux_11 cmd_mux_011(
	.h2f_ARVALID_0(h2f_ARVALID_0),
	.h2f_ARADDR_4(h2f_ARADDR_4),
	.h2f_ARADDR_5(h2f_ARADDR_5),
	.h2f_ARADDR_6(h2f_ARADDR_6),
	.h2f_ARADDR_7(h2f_ARADDR_7),
	.h2f_ARADDR_8(h2f_ARADDR_8),
	.h2f_ARSIZE_0(h2f_ARSIZE_0),
	.h2f_ARSIZE_1(h2f_ARSIZE_1),
	.h2f_ARSIZE_2(h2f_ARSIZE_2),
	.has_pending_responses(\hps_0_h2f_axi_master_rd_limiter|has_pending_responses~q ),
	.saved_grant_1(\cmd_mux_011|saved_grant[1]~q ),
	.last_cycle(\cmd_mux_011|last_cycle~0_combout ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.nxt_in_ready(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.last_channel_11(\hps_0_h2f_axi_master_rd_limiter|last_channel[11]~q ),
	.src_valid(\cmd_mux_011|src_valid~0_combout ),
	.src_payload(\cmd_mux_011|src_payload~0_combout ),
	.src_payload1(\cmd_mux_011|src_payload~1_combout ),
	.src_payload2(\cmd_mux_011|src_payload~2_combout ),
	.clk_clk(clk_clk));

spw_babasu_spw_babasu_mm_interconnect_0_cmd_mux_10 cmd_mux_010(
	.h2f_ARVALID_0(h2f_ARVALID_0),
	.h2f_ARSIZE_0(h2f_ARSIZE_0),
	.h2f_ARSIZE_1(h2f_ARSIZE_1),
	.h2f_ARSIZE_2(h2f_ARSIZE_2),
	.has_pending_responses(\hps_0_h2f_axi_master_rd_limiter|has_pending_responses~q ),
	.saved_grant_1(\cmd_mux_010|saved_grant[1]~q ),
	.Equal10(\router_001|Equal10~0_combout ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.last_channel_10(\hps_0_h2f_axi_master_rd_limiter|last_channel[10]~q ),
	.src_valid(\cmd_mux_010|src_valid~0_combout ),
	.nxt_in_ready(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.src_payload(\cmd_mux_010|src_payload~0_combout ),
	.src_payload1(\cmd_mux_010|src_payload~1_combout ),
	.src_payload2(\cmd_mux_010|src_payload~2_combout ),
	.clk_clk(clk_clk));

spw_babasu_spw_babasu_mm_interconnect_0_rsp_mux_1 rsp_mux_001(
	.read_latency_shift_reg_0(\wr_data_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\wr_data_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_66_0(\wr_data_s1_agent_rsp_fifo|mem[0][66]~q ),
	.read_latency_shift_reg_01(\rd_data_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_01(\rd_data_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_66_01(\rd_data_s1_agent_rsp_fifo|mem[0][66]~q ),
	.read_latency_shift_reg_02(\link_start_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_02(\link_start_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_66_02(\link_start_s1_agent_rsp_fifo|mem[0][66]~q ),
	.read_latency_shift_reg_03(\link_disable_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_03(\link_disable_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_66_03(\link_disable_s1_agent_rsp_fifo|mem[0][66]~q ),
	.read_latency_shift_reg_04(\autostart_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_04(\autostart_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_66_04(\autostart_s1_agent_rsp_fifo|mem[0][66]~q ),
	.mem_66_05(\data_i_s1_agent_rsp_fifo|mem[0][66]~q ),
	.read_latency_shift_reg_05(\tick_in_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_05(\tick_in_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_66_06(\tick_in_s1_agent_rsp_fifo|mem[0][66]~q ),
	.mem_66_07(\time_in_s1_agent_rsp_fifo|mem[0][66]~q ),
	.mem_66_08(\tx_clk_div_s1_agent_rsp_fifo|mem[0][66]~q ),
	.read_latency_shift_reg_06(\spill_enable_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_06(\spill_enable_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_66_09(\spill_enable_s1_agent_rsp_fifo|mem[0][66]~q ),
	.comb(\spill_enable_s1_agent|comb~0_combout ),
	.src1_valid(\rsp_demux_016|src1_valid~0_combout ),
	.mem_130_0(\spill_enable_s1_agent_rsp_fifo|mem[0][130]~q ),
	.last_packet_beat(\spill_enable_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.last_packet_beat1(\spill_enable_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.src_payload(\rsp_mux_001|src_payload~0_combout ),
	.read_latency_shift_reg_07(\tx_full_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_07(\tx_full_s1_agent_rdata_fifo|mem_used[0]~q ),
	.empty(\tx_full_s1_agent_rdata_fifo|empty~combout ),
	.last_packet_beat2(\tx_full_s1_agent|uncompressor|last_packet_beat~3_combout ),
	.mem_130_01(\time_out_s1_agent_rsp_fifo|mem[0][130]~q ),
	.read_latency_shift_reg_08(\time_out_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_08(\time_out_s1_agent_rdata_fifo|mem_used[0]~q ),
	.empty1(\time_out_s1_agent_rdata_fifo|empty~combout ),
	.mem_66_010(\time_out_s1_agent_rsp_fifo|mem[0][66]~q ),
	.mem_used_09(\time_out_s1_agent_rsp_fifo|mem_used[0]~q ),
	.last_packet_beat3(\time_out_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.last_packet_beat4(\time_out_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.mem_130_02(\tick_out_s1_agent_rsp_fifo|mem[0][130]~q ),
	.read_latency_shift_reg_09(\tick_out_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_010(\tick_out_s1_agent_rdata_fifo|mem_used[0]~q ),
	.empty2(\tick_out_s1_agent_rdata_fifo|empty~combout ),
	.mem_66_011(\tick_out_s1_agent_rsp_fifo|mem[0][66]~q ),
	.mem_used_011(\tick_out_s1_agent_rsp_fifo|mem_used[0]~q ),
	.last_packet_beat5(\tick_out_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.last_packet_beat6(\tick_out_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.mem_130_03(\rx_empty_s1_agent_rsp_fifo|mem[0][130]~q ),
	.read_latency_shift_reg_010(\rx_empty_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_012(\rx_empty_s1_agent_rdata_fifo|mem_used[0]~q ),
	.empty3(\rx_empty_s1_agent_rdata_fifo|empty~combout ),
	.mem_66_012(\rx_empty_s1_agent_rsp_fifo|mem[0][66]~q ),
	.mem_used_013(\rx_empty_s1_agent_rsp_fifo|mem_used[0]~q ),
	.last_packet_beat7(\rx_empty_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.last_packet_beat8(\rx_empty_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.mem_130_04(\tx_full_s1_agent_rsp_fifo|mem[0][130]~q ),
	.mem_130_05(\data_o_s1_agent_rsp_fifo|mem[0][130]~q ),
	.read_latency_shift_reg_011(\data_o_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_014(\data_o_s1_agent_rdata_fifo|mem_used[0]~q ),
	.empty4(\data_o_s1_agent_rdata_fifo|empty~combout ),
	.mem_66_013(\data_o_s1_agent_rsp_fifo|mem[0][66]~q ),
	.mem_used_015(\data_o_s1_agent_rsp_fifo|mem_used[0]~q ),
	.last_packet_beat9(\data_o_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.last_packet_beat10(\data_o_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.src_payload_0(\rsp_mux_001|src_payload[0]~6_combout ),
	.comb1(\link_start_s1_agent|comb~0_combout ),
	.src1_valid1(\rsp_demux|src1_valid~0_combout ),
	.mem_130_06(\link_start_s1_agent_rsp_fifo|mem[0][130]~q ),
	.last_packet_beat11(\link_start_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.last_packet_beat12(\link_start_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.comb2(\link_disable_s1_agent|comb~0_combout ),
	.src1_valid2(\rsp_demux_001|src1_valid~0_combout ),
	.mem_130_07(\link_disable_s1_agent_rsp_fifo|mem[0][130]~q ),
	.last_packet_beat13(\link_disable_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.last_packet_beat14(\link_disable_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.comb3(\autostart_s1_agent|comb~0_combout ),
	.src1_valid3(\rsp_demux_002|src1_valid~0_combout ),
	.mem_130_08(\autostart_s1_agent_rsp_fifo|mem[0][130]~q ),
	.last_packet_beat15(\autostart_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.last_packet_beat16(\autostart_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.comb4(\data_i_s1_agent|comb~0_combout ),
	.src1_valid4(\rsp_demux_005|src1_valid~0_combout ),
	.mem_130_09(\data_i_s1_agent_rsp_fifo|mem[0][130]~q ),
	.last_packet_beat17(\data_i_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.last_packet_beat18(\data_i_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.comb5(\wr_data_s1_agent|comb~0_combout ),
	.src1_valid5(\rsp_demux_006|src1_valid~0_combout ),
	.mem_130_010(\wr_data_s1_agent_rsp_fifo|mem[0][130]~q ),
	.last_packet_beat19(\wr_data_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.last_packet_beat20(\wr_data_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.mem_130_011(\currentstate_s1_agent_rsp_fifo|mem[0][130]~q ),
	.read_latency_shift_reg_012(\currentstate_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_016(\currentstate_s1_agent_rdata_fifo|mem_used[0]~q ),
	.empty5(\currentstate_s1_agent_rdata_fifo|empty~combout ),
	.mem_66_014(\currentstate_s1_agent_rsp_fifo|mem[0][66]~q ),
	.mem_used_017(\currentstate_s1_agent_rsp_fifo|mem_used[0]~q ),
	.last_packet_beat21(\currentstate_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.last_packet_beat22(\currentstate_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.src_payload_01(\rsp_mux_001|src_payload[0]~13_combout ),
	.read_latency_shift_reg_013(\flags_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_018(\flags_s1_agent_rdata_fifo|mem_used[0]~q ),
	.empty6(\flags_s1_agent_rdata_fifo|empty~combout ),
	.last_packet_beat23(\flags_s1_agent|uncompressor|last_packet_beat~3_combout ),
	.comb6(\rd_data_s1_agent|comb~0_combout ),
	.src1_valid6(\rsp_demux_009|src1_valid~0_combout ),
	.mem_130_012(\rd_data_s1_agent_rsp_fifo|mem[0][130]~q ),
	.last_packet_beat24(\rd_data_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.last_packet_beat25(\rd_data_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.comb7(\tick_in_s1_agent|comb~0_combout ),
	.src1_valid7(\rsp_demux_013|src1_valid~0_combout ),
	.mem_130_013(\tick_in_s1_agent_rsp_fifo|mem[0][130]~q ),
	.last_packet_beat26(\tick_in_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.last_packet_beat27(\tick_in_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.comb8(\time_in_s1_agent|comb~0_combout ),
	.src1_valid8(\rsp_demux_014|src1_valid~0_combout ),
	.mem_130_014(\time_in_s1_agent_rsp_fifo|mem[0][130]~q ),
	.last_packet_beat28(\time_in_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.last_packet_beat29(\time_in_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.comb9(\tx_clk_div_s1_agent|comb~0_combout ),
	.src1_valid9(\rsp_demux_015|src1_valid~0_combout ),
	.mem_130_015(\tx_clk_div_s1_agent_rsp_fifo|mem[0][130]~q ),
	.last_packet_beat30(\tx_clk_div_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.last_packet_beat31(\tx_clk_div_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.mem_130_016(\flags_s1_agent_rsp_fifo|mem[0][130]~q ),
	.src_payload_02(\rsp_mux_001|src_payload[0]~19_combout ),
	.src_payload_03(src_payload_0),
	.WideOr11(WideOr11),
	.mem_105_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][105]~q ),
	.mem_105_01(\spill_enable_s1_agent_rsp_fifo|mem[0][105]~q ),
	.mem_105_02(\tick_in_s1_agent_rsp_fifo|mem[0][105]~q ),
	.mem_105_03(\time_in_s1_agent_rsp_fifo|mem[0][105]~q ),
	.mem_105_04(\autostart_s1_agent_rsp_fifo|mem[0][105]~q ),
	.mem_105_05(\rd_data_s1_agent_rsp_fifo|mem[0][105]~q ),
	.mem_105_06(\link_start_s1_agent_rsp_fifo|mem[0][105]~q ),
	.mem_105_07(\link_disable_s1_agent_rsp_fifo|mem[0][105]~q ),
	.mem_105_08(\data_i_s1_agent_rsp_fifo|mem[0][105]~q ),
	.mem_105_09(\wr_data_s1_agent_rsp_fifo|mem[0][105]~q ),
	.mem_106_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][106]~q ),
	.mem_106_01(\spill_enable_s1_agent_rsp_fifo|mem[0][106]~q ),
	.mem_106_02(\tick_in_s1_agent_rsp_fifo|mem[0][106]~q ),
	.mem_106_03(\time_in_s1_agent_rsp_fifo|mem[0][106]~q ),
	.mem_106_04(\autostart_s1_agent_rsp_fifo|mem[0][106]~q ),
	.mem_106_05(\rd_data_s1_agent_rsp_fifo|mem[0][106]~q ),
	.mem_106_06(\link_start_s1_agent_rsp_fifo|mem[0][106]~q ),
	.mem_106_07(\link_disable_s1_agent_rsp_fifo|mem[0][106]~q ),
	.mem_106_08(\data_i_s1_agent_rsp_fifo|mem[0][106]~q ),
	.mem_106_09(\wr_data_s1_agent_rsp_fifo|mem[0][106]~q ),
	.mem_107_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][107]~q ),
	.mem_107_01(\spill_enable_s1_agent_rsp_fifo|mem[0][107]~q ),
	.mem_107_02(\tick_in_s1_agent_rsp_fifo|mem[0][107]~q ),
	.mem_107_03(\time_in_s1_agent_rsp_fifo|mem[0][107]~q ),
	.mem_107_04(\autostart_s1_agent_rsp_fifo|mem[0][107]~q ),
	.mem_107_05(\rd_data_s1_agent_rsp_fifo|mem[0][107]~q ),
	.mem_107_06(\link_start_s1_agent_rsp_fifo|mem[0][107]~q ),
	.mem_107_07(\link_disable_s1_agent_rsp_fifo|mem[0][107]~q ),
	.mem_107_08(\data_i_s1_agent_rsp_fifo|mem[0][107]~q ),
	.mem_107_09(\wr_data_s1_agent_rsp_fifo|mem[0][107]~q ),
	.mem_108_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][108]~q ),
	.mem_108_01(\spill_enable_s1_agent_rsp_fifo|mem[0][108]~q ),
	.mem_108_02(\tick_in_s1_agent_rsp_fifo|mem[0][108]~q ),
	.mem_108_03(\time_in_s1_agent_rsp_fifo|mem[0][108]~q ),
	.mem_108_04(\autostart_s1_agent_rsp_fifo|mem[0][108]~q ),
	.mem_108_05(\rd_data_s1_agent_rsp_fifo|mem[0][108]~q ),
	.mem_108_06(\link_start_s1_agent_rsp_fifo|mem[0][108]~q ),
	.mem_108_07(\link_disable_s1_agent_rsp_fifo|mem[0][108]~q ),
	.mem_108_08(\data_i_s1_agent_rsp_fifo|mem[0][108]~q ),
	.mem_108_09(\wr_data_s1_agent_rsp_fifo|mem[0][108]~q ),
	.mem_109_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][109]~q ),
	.mem_109_01(\spill_enable_s1_agent_rsp_fifo|mem[0][109]~q ),
	.mem_109_02(\tick_in_s1_agent_rsp_fifo|mem[0][109]~q ),
	.mem_109_03(\time_in_s1_agent_rsp_fifo|mem[0][109]~q ),
	.mem_109_04(\autostart_s1_agent_rsp_fifo|mem[0][109]~q ),
	.mem_109_05(\rd_data_s1_agent_rsp_fifo|mem[0][109]~q ),
	.mem_109_06(\link_start_s1_agent_rsp_fifo|mem[0][109]~q ),
	.mem_109_07(\link_disable_s1_agent_rsp_fifo|mem[0][109]~q ),
	.mem_109_08(\data_i_s1_agent_rsp_fifo|mem[0][109]~q ),
	.mem_109_09(\wr_data_s1_agent_rsp_fifo|mem[0][109]~q ),
	.mem_110_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][110]~q ),
	.mem_110_01(\spill_enable_s1_agent_rsp_fifo|mem[0][110]~q ),
	.mem_110_02(\tick_in_s1_agent_rsp_fifo|mem[0][110]~q ),
	.mem_110_03(\time_in_s1_agent_rsp_fifo|mem[0][110]~q ),
	.mem_110_04(\autostart_s1_agent_rsp_fifo|mem[0][110]~q ),
	.mem_110_05(\rd_data_s1_agent_rsp_fifo|mem[0][110]~q ),
	.mem_110_06(\link_start_s1_agent_rsp_fifo|mem[0][110]~q ),
	.mem_110_07(\link_disable_s1_agent_rsp_fifo|mem[0][110]~q ),
	.mem_110_08(\data_i_s1_agent_rsp_fifo|mem[0][110]~q ),
	.mem_110_09(\wr_data_s1_agent_rsp_fifo|mem[0][110]~q ),
	.mem_111_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][111]~q ),
	.mem_111_01(\spill_enable_s1_agent_rsp_fifo|mem[0][111]~q ),
	.mem_111_02(\tick_in_s1_agent_rsp_fifo|mem[0][111]~q ),
	.mem_111_03(\time_in_s1_agent_rsp_fifo|mem[0][111]~q ),
	.mem_111_04(\autostart_s1_agent_rsp_fifo|mem[0][111]~q ),
	.mem_111_05(\rd_data_s1_agent_rsp_fifo|mem[0][111]~q ),
	.mem_111_06(\link_start_s1_agent_rsp_fifo|mem[0][111]~q ),
	.mem_111_07(\link_disable_s1_agent_rsp_fifo|mem[0][111]~q ),
	.mem_111_08(\data_i_s1_agent_rsp_fifo|mem[0][111]~q ),
	.mem_111_09(\wr_data_s1_agent_rsp_fifo|mem[0][111]~q ),
	.mem_112_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_112_01(\spill_enable_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_112_02(\tick_in_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_112_03(\time_in_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_112_04(\autostart_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_112_05(\rd_data_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_112_06(\link_start_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_112_07(\link_disable_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_112_08(\data_i_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_112_09(\wr_data_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_113_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][113]~q ),
	.mem_113_01(\spill_enable_s1_agent_rsp_fifo|mem[0][113]~q ),
	.mem_113_02(\tick_in_s1_agent_rsp_fifo|mem[0][113]~q ),
	.mem_113_03(\time_in_s1_agent_rsp_fifo|mem[0][113]~q ),
	.mem_113_04(\autostart_s1_agent_rsp_fifo|mem[0][113]~q ),
	.mem_113_05(\rd_data_s1_agent_rsp_fifo|mem[0][113]~q ),
	.mem_113_06(\link_start_s1_agent_rsp_fifo|mem[0][113]~q ),
	.mem_113_07(\link_disable_s1_agent_rsp_fifo|mem[0][113]~q ),
	.mem_113_08(\data_i_s1_agent_rsp_fifo|mem[0][113]~q ),
	.mem_113_09(\wr_data_s1_agent_rsp_fifo|mem[0][113]~q ),
	.mem_114_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][114]~q ),
	.mem_114_01(\spill_enable_s1_agent_rsp_fifo|mem[0][114]~q ),
	.mem_114_02(\tick_in_s1_agent_rsp_fifo|mem[0][114]~q ),
	.mem_114_03(\time_in_s1_agent_rsp_fifo|mem[0][114]~q ),
	.mem_114_04(\autostart_s1_agent_rsp_fifo|mem[0][114]~q ),
	.mem_114_05(\rd_data_s1_agent_rsp_fifo|mem[0][114]~q ),
	.mem_114_06(\link_start_s1_agent_rsp_fifo|mem[0][114]~q ),
	.mem_114_07(\link_disable_s1_agent_rsp_fifo|mem[0][114]~q ),
	.mem_114_08(\data_i_s1_agent_rsp_fifo|mem[0][114]~q ),
	.mem_114_09(\wr_data_s1_agent_rsp_fifo|mem[0][114]~q ),
	.mem_115_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][115]~q ),
	.mem_115_01(\spill_enable_s1_agent_rsp_fifo|mem[0][115]~q ),
	.mem_115_02(\tick_in_s1_agent_rsp_fifo|mem[0][115]~q ),
	.mem_115_03(\time_in_s1_agent_rsp_fifo|mem[0][115]~q ),
	.mem_115_04(\autostart_s1_agent_rsp_fifo|mem[0][115]~q ),
	.mem_115_05(\rd_data_s1_agent_rsp_fifo|mem[0][115]~q ),
	.mem_115_06(\link_start_s1_agent_rsp_fifo|mem[0][115]~q ),
	.mem_115_07(\link_disable_s1_agent_rsp_fifo|mem[0][115]~q ),
	.mem_115_08(\data_i_s1_agent_rsp_fifo|mem[0][115]~q ),
	.mem_115_09(\wr_data_s1_agent_rsp_fifo|mem[0][115]~q ),
	.mem_116_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][116]~q ),
	.mem_116_01(\spill_enable_s1_agent_rsp_fifo|mem[0][116]~q ),
	.mem_116_02(\tick_in_s1_agent_rsp_fifo|mem[0][116]~q ),
	.mem_116_03(\time_in_s1_agent_rsp_fifo|mem[0][116]~q ),
	.mem_116_04(\autostart_s1_agent_rsp_fifo|mem[0][116]~q ),
	.mem_116_05(\rd_data_s1_agent_rsp_fifo|mem[0][116]~q ),
	.mem_116_06(\link_start_s1_agent_rsp_fifo|mem[0][116]~q ),
	.mem_116_07(\link_disable_s1_agent_rsp_fifo|mem[0][116]~q ),
	.mem_116_08(\data_i_s1_agent_rsp_fifo|mem[0][116]~q ),
	.mem_116_09(\wr_data_s1_agent_rsp_fifo|mem[0][116]~q ),
	.av_readdata_pre_0(\autostart_s1_translator|av_readdata_pre[0]~q ),
	.mem_0_0(\autostart_s1_agent_rdata_fifo|mem[0][0]~q ),
	.av_readdata_pre_01(\tx_clk_div_s1_translator|av_readdata_pre[0]~q ),
	.always4(\tx_clk_div_s1_agent_rdata_fifo|always4~0_combout ),
	.mem_0_01(\tx_clk_div_s1_agent_rdata_fifo|mem[0][0]~q ),
	.av_readdata_pre_02(\currentstate_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_03(\data_o_s1_translator|av_readdata_pre[0]~q ),
	.mem_0_02(\tx_full_s1_agent_rdata_fifo|mem[0][0]~q ),
	.av_readdata_pre_04(\tx_full_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_05(\flags_s1_translator|av_readdata_pre[0]~q ),
	.mem_0_03(\flags_s1_agent_rdata_fifo|mem[0][0]~q ),
	.mem_0_04(\time_out_s1_agent_rdata_fifo|mem[0][0]~q ),
	.av_readdata_pre_06(\time_out_s1_translator|av_readdata_pre[0]~q ),
	.mem_0_05(\data_o_s1_agent_rdata_fifo|mem[0][0]~q ),
	.av_readdata_pre_07(\tick_out_s1_translator|av_readdata_pre[0]~q ),
	.mem_0_06(\tick_out_s1_agent_rdata_fifo|mem[0][0]~q ),
	.av_readdata_pre_08(\rx_empty_s1_translator|av_readdata_pre[0]~q ),
	.mem_0_07(\currentstate_s1_agent_rdata_fifo|mem[0][0]~q ),
	.mem_0_08(\rx_empty_s1_agent_rdata_fifo|mem[0][0]~q ),
	.av_readdata_pre_09(\link_start_s1_translator|av_readdata_pre[0]~q ),
	.mem_0_09(\link_start_s1_agent_rdata_fifo|mem[0][0]~q ),
	.av_readdata_pre_010(\link_disable_s1_translator|av_readdata_pre[0]~q ),
	.mem_0_010(\link_disable_s1_agent_rdata_fifo|mem[0][0]~q ),
	.av_readdata_pre_011(\wr_data_s1_translator|av_readdata_pre[0]~q ),
	.mem_0_011(\wr_data_s1_agent_rdata_fifo|mem[0][0]~q ),
	.av_readdata_pre_012(\rd_data_s1_translator|av_readdata_pre[0]~q ),
	.mem_0_012(\rd_data_s1_agent_rdata_fifo|mem[0][0]~q ),
	.av_readdata_pre_013(\tick_in_s1_translator|av_readdata_pre[0]~q ),
	.mem_0_013(\tick_in_s1_agent_rdata_fifo|mem[0][0]~q ),
	.av_readdata_pre_014(\spill_enable_s1_translator|av_readdata_pre[0]~q ),
	.mem_0_014(\spill_enable_s1_agent_rdata_fifo|mem[0][0]~q ),
	.av_readdata_pre_015(\data_i_s1_translator|av_readdata_pre[0]~q ),
	.always41(\data_i_s1_agent_rdata_fifo|always4~0_combout ),
	.mem_0_015(\data_i_s1_agent_rdata_fifo|mem[0][0]~q ),
	.av_readdata_pre_016(\time_in_s1_translator|av_readdata_pre[0]~q ),
	.always42(\time_in_s1_agent_rdata_fifo|always4~0_combout ),
	.mem_0_016(\time_in_s1_agent_rdata_fifo|mem[0][0]~q ),
	.src_data_0(src_data_0),
	.av_readdata_pre_1(\currentstate_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_11(\data_i_s1_translator|av_readdata_pre[1]~q ),
	.mem_1_0(\data_i_s1_agent_rdata_fifo|mem[0][1]~q ),
	.mem_1_01(\data_o_s1_agent_rdata_fifo|mem[0][1]~q ),
	.mem_1_02(\time_out_s1_agent_rdata_fifo|mem[0][1]~q ),
	.av_readdata_pre_12(\time_out_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_13(\data_o_s1_translator|av_readdata_pre[1]~q ),
	.mem_1_03(\flags_s1_agent_rdata_fifo|mem[0][1]~q ),
	.av_readdata_pre_14(\flags_s1_translator|av_readdata_pre[1]~q ),
	.mem_1_04(\currentstate_s1_agent_rdata_fifo|mem[0][1]~q ),
	.av_readdata_pre_15(\time_in_s1_translator|av_readdata_pre[1]~q ),
	.mem_1_05(\time_in_s1_agent_rdata_fifo|mem[0][1]~q ),
	.av_readdata_pre_16(\tx_clk_div_s1_translator|av_readdata_pre[1]~q ),
	.mem_1_06(\tx_clk_div_s1_agent_rdata_fifo|mem[0][1]~q ),
	.src_payload1(src_payload),
	.av_readdata_pre_2(\currentstate_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_21(\data_i_s1_translator|av_readdata_pre[2]~q ),
	.mem_2_0(\data_i_s1_agent_rdata_fifo|mem[0][2]~q ),
	.mem_2_01(\data_o_s1_agent_rdata_fifo|mem[0][2]~q ),
	.mem_2_02(\time_out_s1_agent_rdata_fifo|mem[0][2]~q ),
	.av_readdata_pre_22(\time_out_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_23(\data_o_s1_translator|av_readdata_pre[2]~q ),
	.mem_2_03(\flags_s1_agent_rdata_fifo|mem[0][2]~q ),
	.av_readdata_pre_24(\flags_s1_translator|av_readdata_pre[2]~q ),
	.mem_2_04(\currentstate_s1_agent_rdata_fifo|mem[0][2]~q ),
	.av_readdata_pre_25(\time_in_s1_translator|av_readdata_pre[2]~q ),
	.mem_2_05(\time_in_s1_agent_rdata_fifo|mem[0][2]~q ),
	.av_readdata_pre_26(\tx_clk_div_s1_translator|av_readdata_pre[2]~q ),
	.mem_2_06(\tx_clk_div_s1_agent_rdata_fifo|mem[0][2]~q ),
	.src_payload2(src_payload1),
	.av_readdata_pre_3(\flags_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_31(\data_i_s1_translator|av_readdata_pre[3]~q ),
	.mem_3_0(\data_i_s1_agent_rdata_fifo|mem[0][3]~q ),
	.mem_3_01(\data_o_s1_agent_rdata_fifo|mem[0][3]~q ),
	.mem_3_02(\time_out_s1_agent_rdata_fifo|mem[0][3]~q ),
	.av_readdata_pre_32(\time_out_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_33(\data_o_s1_translator|av_readdata_pre[3]~q ),
	.mem_3_03(\flags_s1_agent_rdata_fifo|mem[0][3]~q ),
	.av_readdata_pre_34(\time_in_s1_translator|av_readdata_pre[3]~q ),
	.mem_3_04(\time_in_s1_agent_rdata_fifo|mem[0][3]~q ),
	.av_readdata_pre_35(\tx_clk_div_s1_translator|av_readdata_pre[3]~q ),
	.mem_3_05(\tx_clk_div_s1_agent_rdata_fifo|mem[0][3]~q ),
	.src_payload3(src_payload2),
	.av_readdata_pre_4(\flags_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_41(\data_i_s1_translator|av_readdata_pre[4]~q ),
	.mem_4_0(\data_i_s1_agent_rdata_fifo|mem[0][4]~q ),
	.mem_4_01(\data_o_s1_agent_rdata_fifo|mem[0][4]~q ),
	.mem_4_02(\time_out_s1_agent_rdata_fifo|mem[0][4]~q ),
	.av_readdata_pre_42(\time_out_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_43(\data_o_s1_translator|av_readdata_pre[4]~q ),
	.mem_4_03(\flags_s1_agent_rdata_fifo|mem[0][4]~q ),
	.av_readdata_pre_44(\time_in_s1_translator|av_readdata_pre[4]~q ),
	.mem_4_04(\time_in_s1_agent_rdata_fifo|mem[0][4]~q ),
	.av_readdata_pre_45(\tx_clk_div_s1_translator|av_readdata_pre[4]~q ),
	.mem_4_05(\tx_clk_div_s1_agent_rdata_fifo|mem[0][4]~q ),
	.src_payload4(src_payload3),
	.av_readdata_pre_5(\flags_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_51(\data_i_s1_translator|av_readdata_pre[5]~q ),
	.mem_5_0(\data_i_s1_agent_rdata_fifo|mem[0][5]~q ),
	.mem_5_01(\data_o_s1_agent_rdata_fifo|mem[0][5]~q ),
	.mem_5_02(\time_out_s1_agent_rdata_fifo|mem[0][5]~q ),
	.av_readdata_pre_52(\time_out_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_53(\data_o_s1_translator|av_readdata_pre[5]~q ),
	.mem_5_03(\flags_s1_agent_rdata_fifo|mem[0][5]~q ),
	.av_readdata_pre_54(\time_in_s1_translator|av_readdata_pre[5]~q ),
	.mem_5_04(\time_in_s1_agent_rdata_fifo|mem[0][5]~q ),
	.av_readdata_pre_55(\tx_clk_div_s1_translator|av_readdata_pre[5]~q ),
	.mem_5_05(\tx_clk_div_s1_agent_rdata_fifo|mem[0][5]~q ),
	.src_payload5(src_payload4),
	.av_readdata_pre_6(\flags_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_61(\data_i_s1_translator|av_readdata_pre[6]~q ),
	.mem_6_0(\data_i_s1_agent_rdata_fifo|mem[0][6]~q ),
	.mem_6_01(\data_o_s1_agent_rdata_fifo|mem[0][6]~q ),
	.mem_6_02(\time_out_s1_agent_rdata_fifo|mem[0][6]~q ),
	.av_readdata_pre_62(\time_out_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_63(\data_o_s1_translator|av_readdata_pre[6]~q ),
	.mem_6_03(\flags_s1_agent_rdata_fifo|mem[0][6]~q ),
	.av_readdata_pre_64(\time_in_s1_translator|av_readdata_pre[6]~q ),
	.mem_6_04(\time_in_s1_agent_rdata_fifo|mem[0][6]~q ),
	.av_readdata_pre_65(\tx_clk_div_s1_translator|av_readdata_pre[6]~q ),
	.mem_6_05(\tx_clk_div_s1_agent_rdata_fifo|mem[0][6]~q ),
	.src_payload6(src_payload5),
	.av_readdata_pre_7(\flags_s1_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_71(\data_i_s1_translator|av_readdata_pre[7]~q ),
	.mem_7_0(\data_i_s1_agent_rdata_fifo|mem[0][7]~q ),
	.av_readdata_pre_72(\time_in_s1_translator|av_readdata_pre[7]~q ),
	.mem_7_01(\time_in_s1_agent_rdata_fifo|mem[0][7]~q ),
	.mem_7_02(\data_o_s1_agent_rdata_fifo|mem[0][7]~q ),
	.mem_7_03(\time_out_s1_agent_rdata_fifo|mem[0][7]~q ),
	.av_readdata_pre_73(\time_out_s1_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_74(\data_o_s1_translator|av_readdata_pre[7]~q ),
	.mem_7_04(\flags_s1_agent_rdata_fifo|mem[0][7]~q ),
	.src_payload7(src_payload6),
	.av_readdata_pre_8(\data_i_s1_translator|av_readdata_pre[8]~q ),
	.mem_8_0(\data_i_s1_agent_rdata_fifo|mem[0][8]~q ),
	.mem_8_01(\flags_s1_agent_rdata_fifo|mem[0][8]~q ),
	.av_readdata_pre_81(\flags_s1_translator|av_readdata_pre[8]~q ),
	.mem_8_02(\data_o_s1_agent_rdata_fifo|mem[0][8]~q ),
	.av_readdata_pre_82(\data_o_s1_translator|av_readdata_pre[8]~q ),
	.src_payload8(src_payload7),
	.mem_9_0(\flags_s1_agent_rdata_fifo|mem[0][9]~q ),
	.av_readdata_pre_9(\flags_s1_translator|av_readdata_pre[9]~q ),
	.src_payload9(src_payload8),
	.mem_10_0(\flags_s1_agent_rdata_fifo|mem[0][10]~q ),
	.av_readdata_pre_10(\flags_s1_translator|av_readdata_pre[10]~q ),
	.src_payload10(src_payload9),
	.mem_105_010(\time_out_s1_agent_rsp_fifo|mem[0][105]~q ),
	.mem_105_011(\currentstate_s1_agent_rsp_fifo|mem[0][105]~q ),
	.mem_105_012(\flags_s1_agent_rsp_fifo|mem[0][105]~q ),
	.mem_105_013(\tx_full_s1_agent_rsp_fifo|mem[0][105]~q ),
	.mem_105_014(\data_o_s1_agent_rsp_fifo|mem[0][105]~q ),
	.mem_105_015(\rx_empty_s1_agent_rsp_fifo|mem[0][105]~q ),
	.mem_105_016(\tick_out_s1_agent_rsp_fifo|mem[0][105]~q ),
	.src_data_105(src_data_1051),
	.mem_106_010(\time_out_s1_agent_rsp_fifo|mem[0][106]~q ),
	.mem_106_011(\currentstate_s1_agent_rsp_fifo|mem[0][106]~q ),
	.mem_106_012(\flags_s1_agent_rsp_fifo|mem[0][106]~q ),
	.mem_106_013(\tx_full_s1_agent_rsp_fifo|mem[0][106]~q ),
	.mem_106_014(\data_o_s1_agent_rsp_fifo|mem[0][106]~q ),
	.mem_106_015(\rx_empty_s1_agent_rsp_fifo|mem[0][106]~q ),
	.mem_106_016(\tick_out_s1_agent_rsp_fifo|mem[0][106]~q ),
	.src_data_106(src_data_1061),
	.mem_107_010(\time_out_s1_agent_rsp_fifo|mem[0][107]~q ),
	.mem_107_011(\currentstate_s1_agent_rsp_fifo|mem[0][107]~q ),
	.mem_107_012(\flags_s1_agent_rsp_fifo|mem[0][107]~q ),
	.mem_107_013(\tx_full_s1_agent_rsp_fifo|mem[0][107]~q ),
	.mem_107_014(\data_o_s1_agent_rsp_fifo|mem[0][107]~q ),
	.mem_107_015(\rx_empty_s1_agent_rsp_fifo|mem[0][107]~q ),
	.mem_107_016(\tick_out_s1_agent_rsp_fifo|mem[0][107]~q ),
	.src_data_107(src_data_1071),
	.mem_108_010(\time_out_s1_agent_rsp_fifo|mem[0][108]~q ),
	.mem_108_011(\currentstate_s1_agent_rsp_fifo|mem[0][108]~q ),
	.mem_108_012(\flags_s1_agent_rsp_fifo|mem[0][108]~q ),
	.mem_108_013(\tx_full_s1_agent_rsp_fifo|mem[0][108]~q ),
	.mem_108_014(\data_o_s1_agent_rsp_fifo|mem[0][108]~q ),
	.mem_108_015(\rx_empty_s1_agent_rsp_fifo|mem[0][108]~q ),
	.mem_108_016(\tick_out_s1_agent_rsp_fifo|mem[0][108]~q ),
	.src_data_108(src_data_1081),
	.mem_109_010(\time_out_s1_agent_rsp_fifo|mem[0][109]~q ),
	.mem_109_011(\currentstate_s1_agent_rsp_fifo|mem[0][109]~q ),
	.mem_109_012(\flags_s1_agent_rsp_fifo|mem[0][109]~q ),
	.mem_109_013(\tx_full_s1_agent_rsp_fifo|mem[0][109]~q ),
	.mem_109_014(\data_o_s1_agent_rsp_fifo|mem[0][109]~q ),
	.mem_109_015(\rx_empty_s1_agent_rsp_fifo|mem[0][109]~q ),
	.mem_109_016(\tick_out_s1_agent_rsp_fifo|mem[0][109]~q ),
	.src_data_109(src_data_1091),
	.mem_110_010(\time_out_s1_agent_rsp_fifo|mem[0][110]~q ),
	.mem_110_011(\currentstate_s1_agent_rsp_fifo|mem[0][110]~q ),
	.mem_110_012(\flags_s1_agent_rsp_fifo|mem[0][110]~q ),
	.mem_110_013(\tx_full_s1_agent_rsp_fifo|mem[0][110]~q ),
	.mem_110_014(\data_o_s1_agent_rsp_fifo|mem[0][110]~q ),
	.mem_110_015(\rx_empty_s1_agent_rsp_fifo|mem[0][110]~q ),
	.mem_110_016(\tick_out_s1_agent_rsp_fifo|mem[0][110]~q ),
	.src_data_110(src_data_1101),
	.mem_111_010(\time_out_s1_agent_rsp_fifo|mem[0][111]~q ),
	.mem_111_011(\currentstate_s1_agent_rsp_fifo|mem[0][111]~q ),
	.mem_111_012(\flags_s1_agent_rsp_fifo|mem[0][111]~q ),
	.mem_111_013(\tx_full_s1_agent_rsp_fifo|mem[0][111]~q ),
	.mem_111_014(\data_o_s1_agent_rsp_fifo|mem[0][111]~q ),
	.mem_111_015(\rx_empty_s1_agent_rsp_fifo|mem[0][111]~q ),
	.mem_111_016(\tick_out_s1_agent_rsp_fifo|mem[0][111]~q ),
	.src_data_111(src_data_1111),
	.mem_112_010(\time_out_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_112_011(\currentstate_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_112_012(\flags_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_112_013(\tx_full_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_112_014(\data_o_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_112_015(\rx_empty_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_112_016(\tick_out_s1_agent_rsp_fifo|mem[0][112]~q ),
	.src_data_112(src_data_1121),
	.mem_113_010(\time_out_s1_agent_rsp_fifo|mem[0][113]~q ),
	.mem_113_011(\currentstate_s1_agent_rsp_fifo|mem[0][113]~q ),
	.mem_113_012(\flags_s1_agent_rsp_fifo|mem[0][113]~q ),
	.mem_113_013(\tx_full_s1_agent_rsp_fifo|mem[0][113]~q ),
	.mem_113_014(\data_o_s1_agent_rsp_fifo|mem[0][113]~q ),
	.mem_113_015(\rx_empty_s1_agent_rsp_fifo|mem[0][113]~q ),
	.mem_113_016(\tick_out_s1_agent_rsp_fifo|mem[0][113]~q ),
	.src_data_113(src_data_1131),
	.mem_114_010(\time_out_s1_agent_rsp_fifo|mem[0][114]~q ),
	.mem_114_011(\currentstate_s1_agent_rsp_fifo|mem[0][114]~q ),
	.mem_114_012(\flags_s1_agent_rsp_fifo|mem[0][114]~q ),
	.mem_114_013(\tx_full_s1_agent_rsp_fifo|mem[0][114]~q ),
	.mem_114_014(\data_o_s1_agent_rsp_fifo|mem[0][114]~q ),
	.mem_114_015(\rx_empty_s1_agent_rsp_fifo|mem[0][114]~q ),
	.mem_114_016(\tick_out_s1_agent_rsp_fifo|mem[0][114]~q ),
	.src_data_114(src_data_1141),
	.mem_115_010(\time_out_s1_agent_rsp_fifo|mem[0][115]~q ),
	.mem_115_011(\currentstate_s1_agent_rsp_fifo|mem[0][115]~q ),
	.mem_115_012(\flags_s1_agent_rsp_fifo|mem[0][115]~q ),
	.mem_115_013(\tx_full_s1_agent_rsp_fifo|mem[0][115]~q ),
	.mem_115_014(\data_o_s1_agent_rsp_fifo|mem[0][115]~q ),
	.mem_115_015(\rx_empty_s1_agent_rsp_fifo|mem[0][115]~q ),
	.mem_115_016(\tick_out_s1_agent_rsp_fifo|mem[0][115]~q ),
	.src_data_115(src_data_1151),
	.mem_116_010(\time_out_s1_agent_rsp_fifo|mem[0][116]~q ),
	.mem_116_011(\currentstate_s1_agent_rsp_fifo|mem[0][116]~q ),
	.mem_116_012(\flags_s1_agent_rsp_fifo|mem[0][116]~q ),
	.mem_116_013(\tx_full_s1_agent_rsp_fifo|mem[0][116]~q ),
	.mem_116_014(\data_o_s1_agent_rsp_fifo|mem[0][116]~q ),
	.mem_116_015(\rx_empty_s1_agent_rsp_fifo|mem[0][116]~q ),
	.mem_116_016(\tick_out_s1_agent_rsp_fifo|mem[0][116]~q ),
	.src_data_116(src_data_1161));

spw_babasu_spw_babasu_mm_interconnect_0_rsp_mux rsp_mux(
	.mem_66_0(\wr_data_s1_agent_rsp_fifo|mem[0][66]~q ),
	.src0_valid(\rsp_demux_006|src0_valid~combout ),
	.mem_66_01(\rd_data_s1_agent_rsp_fifo|mem[0][66]~q ),
	.src0_valid1(\rsp_demux_009|src0_valid~combout ),
	.mem_66_02(\link_start_s1_agent_rsp_fifo|mem[0][66]~q ),
	.src0_valid2(\rsp_demux|src0_valid~combout ),
	.mem_66_03(\link_disable_s1_agent_rsp_fifo|mem[0][66]~q ),
	.src0_valid3(\rsp_demux_001|src0_valid~combout ),
	.mem_66_04(\autostart_s1_agent_rsp_fifo|mem[0][66]~q ),
	.src0_valid4(\rsp_demux_002|src0_valid~combout ),
	.mem_66_05(\data_i_s1_agent_rsp_fifo|mem[0][66]~q ),
	.src0_valid5(\rsp_demux_005|src0_valid~combout ),
	.src0_valid6(\rsp_demux_013|src0_valid~combout ),
	.src0_valid7(\rsp_demux_014|src0_valid~combout ),
	.mem_66_06(\tx_clk_div_s1_agent_rsp_fifo|mem[0][66]~q ),
	.src0_valid8(\rsp_demux_015|src0_valid~combout ),
	.mem_66_07(\spill_enable_s1_agent_rsp_fifo|mem[0][66]~q ),
	.src0_valid9(\rsp_demux_016|src0_valid~combout ),
	.WideOr11(WideOr1),
	.comb(\spill_enable_s1_agent|comb~0_combout ),
	.mem_130_0(\spill_enable_s1_agent_rsp_fifo|mem[0][130]~q ),
	.last_packet_beat(\spill_enable_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.last_packet_beat1(\spill_enable_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.comb1(\link_start_s1_agent|comb~0_combout ),
	.mem_130_01(\link_start_s1_agent_rsp_fifo|mem[0][130]~q ),
	.last_packet_beat2(\link_start_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.last_packet_beat3(\link_start_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.comb2(\link_disable_s1_agent|comb~0_combout ),
	.mem_130_02(\link_disable_s1_agent_rsp_fifo|mem[0][130]~q ),
	.last_packet_beat4(\link_disable_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.last_packet_beat5(\link_disable_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.comb3(\autostart_s1_agent|comb~0_combout ),
	.mem_130_03(\autostart_s1_agent_rsp_fifo|mem[0][130]~q ),
	.last_packet_beat6(\autostart_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.last_packet_beat7(\autostart_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.comb4(\data_i_s1_agent|comb~0_combout ),
	.mem_130_04(\data_i_s1_agent_rsp_fifo|mem[0][130]~q ),
	.last_packet_beat8(\data_i_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.last_packet_beat9(\data_i_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.comb5(\wr_data_s1_agent|comb~0_combout ),
	.mem_130_05(\wr_data_s1_agent_rsp_fifo|mem[0][130]~q ),
	.last_packet_beat10(\wr_data_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.last_packet_beat11(\wr_data_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.comb6(\rd_data_s1_agent|comb~0_combout ),
	.mem_130_06(\rd_data_s1_agent_rsp_fifo|mem[0][130]~q ),
	.last_packet_beat12(\rd_data_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.last_packet_beat13(\rd_data_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.mem_130_07(\tick_in_s1_agent_rsp_fifo|mem[0][130]~q ),
	.mem_130_08(\time_in_s1_agent_rsp_fifo|mem[0][130]~q ),
	.comb7(\tx_clk_div_s1_agent|comb~0_combout ),
	.mem_130_09(\tx_clk_div_s1_agent_rsp_fifo|mem[0][130]~q ),
	.last_packet_beat14(\tx_clk_div_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.last_packet_beat15(\tx_clk_div_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.mem_105_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][105]~q ),
	.mem_105_01(\spill_enable_s1_agent_rsp_fifo|mem[0][105]~q ),
	.mem_105_02(\tick_in_s1_agent_rsp_fifo|mem[0][105]~q ),
	.mem_105_03(\time_in_s1_agent_rsp_fifo|mem[0][105]~q ),
	.mem_105_04(\autostart_s1_agent_rsp_fifo|mem[0][105]~q ),
	.mem_105_05(\rd_data_s1_agent_rsp_fifo|mem[0][105]~q ),
	.mem_105_06(\link_start_s1_agent_rsp_fifo|mem[0][105]~q ),
	.mem_105_07(\link_disable_s1_agent_rsp_fifo|mem[0][105]~q ),
	.mem_105_08(\data_i_s1_agent_rsp_fifo|mem[0][105]~q ),
	.mem_105_09(\wr_data_s1_agent_rsp_fifo|mem[0][105]~q ),
	.src_data_105(src_data_105),
	.mem_106_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][106]~q ),
	.mem_106_01(\spill_enable_s1_agent_rsp_fifo|mem[0][106]~q ),
	.mem_106_02(\tick_in_s1_agent_rsp_fifo|mem[0][106]~q ),
	.mem_106_03(\time_in_s1_agent_rsp_fifo|mem[0][106]~q ),
	.mem_106_04(\autostart_s1_agent_rsp_fifo|mem[0][106]~q ),
	.mem_106_05(\rd_data_s1_agent_rsp_fifo|mem[0][106]~q ),
	.mem_106_06(\link_start_s1_agent_rsp_fifo|mem[0][106]~q ),
	.mem_106_07(\link_disable_s1_agent_rsp_fifo|mem[0][106]~q ),
	.mem_106_08(\data_i_s1_agent_rsp_fifo|mem[0][106]~q ),
	.mem_106_09(\wr_data_s1_agent_rsp_fifo|mem[0][106]~q ),
	.src_data_106(src_data_106),
	.mem_107_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][107]~q ),
	.mem_107_01(\spill_enable_s1_agent_rsp_fifo|mem[0][107]~q ),
	.mem_107_02(\tick_in_s1_agent_rsp_fifo|mem[0][107]~q ),
	.mem_107_03(\time_in_s1_agent_rsp_fifo|mem[0][107]~q ),
	.mem_107_04(\autostart_s1_agent_rsp_fifo|mem[0][107]~q ),
	.mem_107_05(\rd_data_s1_agent_rsp_fifo|mem[0][107]~q ),
	.mem_107_06(\link_start_s1_agent_rsp_fifo|mem[0][107]~q ),
	.mem_107_07(\link_disable_s1_agent_rsp_fifo|mem[0][107]~q ),
	.mem_107_08(\data_i_s1_agent_rsp_fifo|mem[0][107]~q ),
	.mem_107_09(\wr_data_s1_agent_rsp_fifo|mem[0][107]~q ),
	.src_data_107(src_data_107),
	.mem_108_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][108]~q ),
	.mem_108_01(\spill_enable_s1_agent_rsp_fifo|mem[0][108]~q ),
	.mem_108_02(\tick_in_s1_agent_rsp_fifo|mem[0][108]~q ),
	.mem_108_03(\time_in_s1_agent_rsp_fifo|mem[0][108]~q ),
	.mem_108_04(\autostart_s1_agent_rsp_fifo|mem[0][108]~q ),
	.mem_108_05(\rd_data_s1_agent_rsp_fifo|mem[0][108]~q ),
	.mem_108_06(\link_start_s1_agent_rsp_fifo|mem[0][108]~q ),
	.mem_108_07(\link_disable_s1_agent_rsp_fifo|mem[0][108]~q ),
	.mem_108_08(\data_i_s1_agent_rsp_fifo|mem[0][108]~q ),
	.mem_108_09(\wr_data_s1_agent_rsp_fifo|mem[0][108]~q ),
	.src_data_108(src_data_108),
	.mem_109_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][109]~q ),
	.mem_109_01(\spill_enable_s1_agent_rsp_fifo|mem[0][109]~q ),
	.mem_109_02(\tick_in_s1_agent_rsp_fifo|mem[0][109]~q ),
	.mem_109_03(\time_in_s1_agent_rsp_fifo|mem[0][109]~q ),
	.mem_109_04(\autostart_s1_agent_rsp_fifo|mem[0][109]~q ),
	.mem_109_05(\rd_data_s1_agent_rsp_fifo|mem[0][109]~q ),
	.mem_109_06(\link_start_s1_agent_rsp_fifo|mem[0][109]~q ),
	.mem_109_07(\link_disable_s1_agent_rsp_fifo|mem[0][109]~q ),
	.mem_109_08(\data_i_s1_agent_rsp_fifo|mem[0][109]~q ),
	.mem_109_09(\wr_data_s1_agent_rsp_fifo|mem[0][109]~q ),
	.src_data_109(src_data_109),
	.mem_110_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][110]~q ),
	.mem_110_01(\spill_enable_s1_agent_rsp_fifo|mem[0][110]~q ),
	.mem_110_02(\tick_in_s1_agent_rsp_fifo|mem[0][110]~q ),
	.mem_110_03(\time_in_s1_agent_rsp_fifo|mem[0][110]~q ),
	.mem_110_04(\autostart_s1_agent_rsp_fifo|mem[0][110]~q ),
	.mem_110_05(\rd_data_s1_agent_rsp_fifo|mem[0][110]~q ),
	.mem_110_06(\link_start_s1_agent_rsp_fifo|mem[0][110]~q ),
	.mem_110_07(\link_disable_s1_agent_rsp_fifo|mem[0][110]~q ),
	.mem_110_08(\data_i_s1_agent_rsp_fifo|mem[0][110]~q ),
	.mem_110_09(\wr_data_s1_agent_rsp_fifo|mem[0][110]~q ),
	.src_data_110(src_data_110),
	.mem_111_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][111]~q ),
	.mem_111_01(\spill_enable_s1_agent_rsp_fifo|mem[0][111]~q ),
	.mem_111_02(\tick_in_s1_agent_rsp_fifo|mem[0][111]~q ),
	.mem_111_03(\time_in_s1_agent_rsp_fifo|mem[0][111]~q ),
	.mem_111_04(\autostart_s1_agent_rsp_fifo|mem[0][111]~q ),
	.mem_111_05(\rd_data_s1_agent_rsp_fifo|mem[0][111]~q ),
	.mem_111_06(\link_start_s1_agent_rsp_fifo|mem[0][111]~q ),
	.mem_111_07(\link_disable_s1_agent_rsp_fifo|mem[0][111]~q ),
	.mem_111_08(\data_i_s1_agent_rsp_fifo|mem[0][111]~q ),
	.mem_111_09(\wr_data_s1_agent_rsp_fifo|mem[0][111]~q ),
	.src_data_111(src_data_111),
	.mem_112_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_112_01(\spill_enable_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_112_02(\tick_in_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_112_03(\time_in_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_112_04(\autostart_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_112_05(\rd_data_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_112_06(\link_start_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_112_07(\link_disable_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_112_08(\data_i_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_112_09(\wr_data_s1_agent_rsp_fifo|mem[0][112]~q ),
	.src_data_112(src_data_112),
	.mem_113_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][113]~q ),
	.mem_113_01(\spill_enable_s1_agent_rsp_fifo|mem[0][113]~q ),
	.mem_113_02(\tick_in_s1_agent_rsp_fifo|mem[0][113]~q ),
	.mem_113_03(\time_in_s1_agent_rsp_fifo|mem[0][113]~q ),
	.mem_113_04(\autostart_s1_agent_rsp_fifo|mem[0][113]~q ),
	.mem_113_05(\rd_data_s1_agent_rsp_fifo|mem[0][113]~q ),
	.mem_113_06(\link_start_s1_agent_rsp_fifo|mem[0][113]~q ),
	.mem_113_07(\link_disable_s1_agent_rsp_fifo|mem[0][113]~q ),
	.mem_113_08(\data_i_s1_agent_rsp_fifo|mem[0][113]~q ),
	.mem_113_09(\wr_data_s1_agent_rsp_fifo|mem[0][113]~q ),
	.src_data_113(src_data_113),
	.mem_114_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][114]~q ),
	.mem_114_01(\spill_enable_s1_agent_rsp_fifo|mem[0][114]~q ),
	.mem_114_02(\tick_in_s1_agent_rsp_fifo|mem[0][114]~q ),
	.mem_114_03(\time_in_s1_agent_rsp_fifo|mem[0][114]~q ),
	.mem_114_04(\autostart_s1_agent_rsp_fifo|mem[0][114]~q ),
	.mem_114_05(\rd_data_s1_agent_rsp_fifo|mem[0][114]~q ),
	.mem_114_06(\link_start_s1_agent_rsp_fifo|mem[0][114]~q ),
	.mem_114_07(\link_disable_s1_agent_rsp_fifo|mem[0][114]~q ),
	.mem_114_08(\data_i_s1_agent_rsp_fifo|mem[0][114]~q ),
	.mem_114_09(\wr_data_s1_agent_rsp_fifo|mem[0][114]~q ),
	.src_data_114(src_data_114),
	.mem_115_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][115]~q ),
	.mem_115_01(\spill_enable_s1_agent_rsp_fifo|mem[0][115]~q ),
	.mem_115_02(\tick_in_s1_agent_rsp_fifo|mem[0][115]~q ),
	.mem_115_03(\time_in_s1_agent_rsp_fifo|mem[0][115]~q ),
	.mem_115_04(\autostart_s1_agent_rsp_fifo|mem[0][115]~q ),
	.mem_115_05(\rd_data_s1_agent_rsp_fifo|mem[0][115]~q ),
	.mem_115_06(\link_start_s1_agent_rsp_fifo|mem[0][115]~q ),
	.mem_115_07(\link_disable_s1_agent_rsp_fifo|mem[0][115]~q ),
	.mem_115_08(\data_i_s1_agent_rsp_fifo|mem[0][115]~q ),
	.mem_115_09(\wr_data_s1_agent_rsp_fifo|mem[0][115]~q ),
	.src_data_115(src_data_115),
	.mem_116_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][116]~q ),
	.mem_116_01(\spill_enable_s1_agent_rsp_fifo|mem[0][116]~q ),
	.mem_116_02(\tick_in_s1_agent_rsp_fifo|mem[0][116]~q ),
	.mem_116_03(\time_in_s1_agent_rsp_fifo|mem[0][116]~q ),
	.mem_116_04(\autostart_s1_agent_rsp_fifo|mem[0][116]~q ),
	.mem_116_05(\rd_data_s1_agent_rsp_fifo|mem[0][116]~q ),
	.mem_116_06(\link_start_s1_agent_rsp_fifo|mem[0][116]~q ),
	.mem_116_07(\link_disable_s1_agent_rsp_fifo|mem[0][116]~q ),
	.mem_116_08(\data_i_s1_agent_rsp_fifo|mem[0][116]~q ),
	.mem_116_09(\wr_data_s1_agent_rsp_fifo|mem[0][116]~q ),
	.src_data_116(src_data_116),
	.last_packet_beat16(\tick_in_s1_agent|uncompressor|last_packet_beat~2_combout ),
	.last_packet_beat17(\time_in_s1_agent|uncompressor|last_packet_beat~2_combout ),
	.src_payload(\rsp_mux|src_payload~0_combout ),
	.src_payload1(\rsp_mux|src_payload~1_combout ),
	.src_payload_0(\rsp_mux|src_payload[0]~8_combout ),
	.src_payload_01(\rsp_mux|src_payload[0]~9_combout ));

spw_babasu_spw_babasu_mm_interconnect_0_rsp_demux_16 rsp_demux_016(
	.h2f_BREADY_0(h2f_BREADY_0),
	.h2f_RREADY_0(h2f_RREADY_0),
	.read_latency_shift_reg_0(\spill_enable_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\spill_enable_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_129_0(\spill_enable_s1_agent_rsp_fifo|mem[0][129]~q ),
	.mem_used_01(\spill_enable_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_68_0(\spill_enable_s1_agent_rsp_fifo|mem[0][68]~q ),
	.mem_66_0(\spill_enable_s1_agent_rsp_fifo|mem[0][66]~q ),
	.src0_valid1(\rsp_demux_016|src0_valid~combout ),
	.src1_valid(\rsp_demux_016|src1_valid~0_combout ),
	.WideOr0(\rsp_demux_016|WideOr0~0_combout ));

spw_babasu_spw_babasu_mm_interconnect_0_rsp_demux_15 rsp_demux_015(
	.h2f_BREADY_0(h2f_BREADY_0),
	.h2f_RREADY_0(h2f_RREADY_0),
	.read_latency_shift_reg_0(\tx_clk_div_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\tx_clk_div_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_129_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][129]~q ),
	.mem_used_01(\tx_clk_div_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_68_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][68]~q ),
	.mem_66_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][66]~q ),
	.src0_valid1(\rsp_demux_015|src0_valid~combout ),
	.src1_valid(\rsp_demux_015|src1_valid~0_combout ),
	.WideOr0(\rsp_demux_015|WideOr0~0_combout ));

spw_babasu_spw_babasu_mm_interconnect_0_rsp_demux_14 rsp_demux_014(
	.h2f_BREADY_0(h2f_BREADY_0),
	.h2f_RREADY_0(h2f_RREADY_0),
	.read_latency_shift_reg_0(\time_in_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\time_in_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_129_0(\time_in_s1_agent_rsp_fifo|mem[0][129]~q ),
	.mem_used_01(\time_in_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_68_0(\time_in_s1_agent_rsp_fifo|mem[0][68]~q ),
	.mem_66_0(\time_in_s1_agent_rsp_fifo|mem[0][66]~q ),
	.src0_valid1(\rsp_demux_014|src0_valid~combout ),
	.src1_valid(\rsp_demux_014|src1_valid~0_combout ),
	.WideOr0(\rsp_demux_014|WideOr0~0_combout ));

spw_babasu_spw_babasu_mm_interconnect_0_rsp_demux_13 rsp_demux_013(
	.h2f_BREADY_0(h2f_BREADY_0),
	.h2f_RREADY_0(h2f_RREADY_0),
	.read_latency_shift_reg_0(\tick_in_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\tick_in_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_129_0(\tick_in_s1_agent_rsp_fifo|mem[0][129]~q ),
	.mem_used_01(\tick_in_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_68_0(\tick_in_s1_agent_rsp_fifo|mem[0][68]~q ),
	.mem_66_0(\tick_in_s1_agent_rsp_fifo|mem[0][66]~q ),
	.src0_valid1(\rsp_demux_013|src0_valid~combout ),
	.src1_valid(\rsp_demux_013|src1_valid~0_combout ),
	.WideOr0(\rsp_demux_013|WideOr0~0_combout ));

spw_babasu_spw_babasu_mm_interconnect_0_rsp_demux_9 rsp_demux_009(
	.h2f_BREADY_0(h2f_BREADY_0),
	.h2f_RREADY_0(h2f_RREADY_0),
	.read_latency_shift_reg_0(\rd_data_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\rd_data_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_129_0(\rd_data_s1_agent_rsp_fifo|mem[0][129]~q ),
	.mem_used_01(\rd_data_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_68_0(\rd_data_s1_agent_rsp_fifo|mem[0][68]~q ),
	.mem_66_0(\rd_data_s1_agent_rsp_fifo|mem[0][66]~q ),
	.src0_valid1(\rsp_demux_009|src0_valid~combout ),
	.src1_valid(\rsp_demux_009|src1_valid~0_combout ),
	.WideOr0(\rsp_demux_009|WideOr0~0_combout ));

spw_babasu_spw_babasu_mm_interconnect_0_rsp_demux_6 rsp_demux_006(
	.h2f_BREADY_0(h2f_BREADY_0),
	.h2f_RREADY_0(h2f_RREADY_0),
	.read_latency_shift_reg_0(\wr_data_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\wr_data_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_129_0(\wr_data_s1_agent_rsp_fifo|mem[0][129]~q ),
	.mem_used_01(\wr_data_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_68_0(\wr_data_s1_agent_rsp_fifo|mem[0][68]~q ),
	.mem_66_0(\wr_data_s1_agent_rsp_fifo|mem[0][66]~q ),
	.src0_valid1(\rsp_demux_006|src0_valid~combout ),
	.src1_valid(\rsp_demux_006|src1_valid~0_combout ),
	.WideOr0(\rsp_demux_006|WideOr0~0_combout ));

spw_babasu_altera_merlin_burst_adapter_3 data_o_s1_burst_adapter(
	.h2f_ARADDR_0(h2f_ARADDR_0),
	.h2f_ARADDR_1(h2f_ARADDR_1),
	.h2f_ARADDR_2(h2f_ARADDR_2),
	.h2f_ARADDR_3(h2f_ARADDR_3),
	.h2f_ARBURST_0(h2f_ARBURST_0),
	.h2f_ARBURST_1(h2f_ARBURST_1),
	.h2f_ARID_0(h2f_ARID_0),
	.h2f_ARID_1(h2f_ARID_1),
	.h2f_ARID_2(h2f_ARID_2),
	.h2f_ARID_3(h2f_ARID_3),
	.h2f_ARID_4(h2f_ARID_4),
	.h2f_ARID_5(h2f_ARID_5),
	.h2f_ARID_6(h2f_ARID_6),
	.h2f_ARID_7(h2f_ARID_7),
	.h2f_ARID_8(h2f_ARID_8),
	.h2f_ARID_9(h2f_ARID_9),
	.h2f_ARID_10(h2f_ARID_10),
	.h2f_ARID_11(h2f_ARID_11),
	.h2f_ARLEN_0(h2f_ARLEN_0),
	.Add5(\hps_0_h2f_axi_master_agent|Add5~1_sumout ),
	.Add51(\hps_0_h2f_axi_master_agent|Add5~5_sumout ),
	.saved_grant_1(\cmd_mux_008|saved_grant[1]~q ),
	.stateST_COMP_TRANS(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.mem_used_1(\data_o_s1_agent_rsp_fifo|mem_used[1]~q ),
	.in_data_reg_69(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.in_narrow_reg(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.cp_ready(\data_o_s1_agent|cp_ready~0_combout ),
	.cp_ready1(\data_o_s1_agent|cp_ready~1_combout ),
	.nxt_out_eop(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.in_ready_hold(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.out_valid_reg(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.stateST_UNCOMP_WR_SUBBURST(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.nxt_in_ready(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.nxt_in_ready1(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.src_valid(\cmd_mux_008|src_valid~0_combout ),
	.Decoder1(\hps_0_h2f_axi_master_agent|Decoder1~0_combout ),
	.out_byte_cnt_reg_2(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.Add2(\hps_0_h2f_axi_master_agent|Add2~0_combout ),
	.Add21(\hps_0_h2f_axi_master_agent|Add2~1_combout ),
	.Add22(\hps_0_h2f_axi_master_agent|Add2~2_combout ),
	.Add23(\hps_0_h2f_axi_master_agent|Add2~3_combout ),
	.cp_ready2(\data_o_s1_agent|cp_ready~2_combout ),
	.out_uncomp_byte_cnt_reg_6(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.out_uncomp_byte_cnt_reg_5(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_4(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_3(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.in_data_reg_105(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ),
	.in_data_reg_106(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ),
	.in_data_reg_107(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ),
	.in_data_reg_108(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ),
	.in_data_reg_109(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ),
	.in_data_reg_110(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ),
	.in_data_reg_111(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ),
	.in_data_reg_112(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ),
	.in_data_reg_113(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ),
	.in_data_reg_114(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ),
	.in_data_reg_115(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ),
	.in_data_reg_116(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ),
	.Selector10(\hps_0_h2f_axi_master_agent|Selector10~0_combout ),
	.Selector101(\hps_0_h2f_axi_master_agent|Selector10~1_combout ),
	.Selector11(\hps_0_h2f_axi_master_agent|Selector11~1_combout ),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_311),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_211),
	.Selector12(\hps_0_h2f_axi_master_agent|Selector12~0_combout ),
	.src_payload(\cmd_mux_008|src_payload~0_combout ),
	.src_payload1(\cmd_mux_008|src_payload~1_combout ),
	.src_payload2(\cmd_mux_008|src_payload~2_combout ),
	.Selector13(\hps_0_h2f_axi_master_agent|Selector13~1_combout ),
	.nxt_out_burstwrap_1(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_burstwrap[1]~0_combout ),
	.nxt_addr_2(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_addr[2]~2_combout ),
	.clk_clk(clk_clk));

spw_babasu_altera_merlin_burst_adapter_15 tx_full_s1_burst_adapter(
	.h2f_ARADDR_0(h2f_ARADDR_0),
	.h2f_ARADDR_1(h2f_ARADDR_1),
	.h2f_ARADDR_2(h2f_ARADDR_2),
	.h2f_ARADDR_3(h2f_ARADDR_3),
	.h2f_ARBURST_0(h2f_ARBURST_0),
	.h2f_ARBURST_1(h2f_ARBURST_1),
	.h2f_ARID_0(h2f_ARID_0),
	.h2f_ARID_1(h2f_ARID_1),
	.h2f_ARID_2(h2f_ARID_2),
	.h2f_ARID_3(h2f_ARID_3),
	.h2f_ARID_4(h2f_ARID_4),
	.h2f_ARID_5(h2f_ARID_5),
	.h2f_ARID_6(h2f_ARID_6),
	.h2f_ARID_7(h2f_ARID_7),
	.h2f_ARID_8(h2f_ARID_8),
	.h2f_ARID_9(h2f_ARID_9),
	.h2f_ARID_10(h2f_ARID_10),
	.h2f_ARID_11(h2f_ARID_11),
	.h2f_ARLEN_0(h2f_ARLEN_0),
	.Add5(\hps_0_h2f_axi_master_agent|Add5~1_sumout ),
	.Add51(\hps_0_h2f_axi_master_agent|Add5~5_sumout ),
	.in_ready_hold(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.in_data_reg_69(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.stateST_COMP_TRANS(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.mem_used_1(\tx_full_s1_agent_rsp_fifo|mem_used[1]~q ),
	.in_narrow_reg(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.cp_ready(\tx_full_s1_agent|cp_ready~0_combout ),
	.nxt_in_ready(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.out_valid_reg(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.stateST_UNCOMP_WR_SUBBURST(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.nxt_in_ready1(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.saved_grant_1(\cmd_mux_007|saved_grant[1]~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.Decoder1(\hps_0_h2f_axi_master_agent|Decoder1~0_combout ),
	.Add2(\hps_0_h2f_axi_master_agent|Add2~0_combout ),
	.Add21(\hps_0_h2f_axi_master_agent|Add2~1_combout ),
	.Add22(\hps_0_h2f_axi_master_agent|Add2~2_combout ),
	.Add23(\hps_0_h2f_axi_master_agent|Add2~3_combout ),
	.nxt_in_ready2(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ),
	.src_valid(\cmd_mux_007|src_valid~0_combout ),
	.nxt_out_eop(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.out_byte_cnt_reg_2(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.cp_ready1(\tx_full_s1_agent|cp_ready~1_combout ),
	.out_uncomp_byte_cnt_reg_3(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_6(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.out_uncomp_byte_cnt_reg_5(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_4(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.in_data_reg_105(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ),
	.in_data_reg_106(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ),
	.in_data_reg_107(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ),
	.in_data_reg_108(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ),
	.in_data_reg_109(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ),
	.in_data_reg_110(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ),
	.in_data_reg_111(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ),
	.in_data_reg_112(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ),
	.in_data_reg_113(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ),
	.in_data_reg_114(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ),
	.in_data_reg_115(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ),
	.in_data_reg_116(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ),
	.Selector10(\hps_0_h2f_axi_master_agent|Selector10~0_combout ),
	.Selector101(\hps_0_h2f_axi_master_agent|Selector10~1_combout ),
	.Selector11(\hps_0_h2f_axi_master_agent|Selector11~1_combout ),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_312),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_212),
	.Selector12(\hps_0_h2f_axi_master_agent|Selector12~0_combout ),
	.src_payload(\cmd_mux_007|src_payload~0_combout ),
	.src_payload1(\cmd_mux_007|src_payload~1_combout ),
	.src_payload2(\cmd_mux_007|src_payload~2_combout ),
	.Selector13(\hps_0_h2f_axi_master_agent|Selector13~1_combout ),
	.nxt_out_burstwrap_1(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_burstwrap[1]~0_combout ),
	.nxt_addr_2(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_addr[2]~2_combout ),
	.clk_clk(clk_clk));

spw_babasu_altera_merlin_burst_adapter_16 wr_data_s1_burst_adapter(
	.h2f_ARADDR_0(h2f_ARADDR_0),
	.h2f_ARADDR_1(h2f_ARADDR_1),
	.h2f_ARADDR_2(h2f_ARADDR_2),
	.h2f_ARADDR_3(h2f_ARADDR_3),
	.h2f_ARLEN_0(h2f_ARLEN_0),
	.nxt_in_ready(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.in_ready_hold(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.stateST_COMP_TRANS(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.out_valid_reg(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.in_narrow_reg(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.in_byteen_reg_3(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ),
	.in_byteen_reg_2(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ),
	.in_byteen_reg_1(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ),
	.in_byteen_reg_0(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ),
	.in_data_reg_68(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ),
	.cp_ready(\wr_data_s1_agent|cp_ready~0_combout ),
	.stateST_UNCOMP_WR_SUBBURST(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.nxt_in_ready1(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.saved_grant_1(\cmd_mux_006|saved_grant[1]~q ),
	.Equal5(\router|Equal5~0_combout ),
	.saved_grant_0(\cmd_mux_006|saved_grant[0]~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.in_data_reg_0(in_data_reg_09),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_39),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_29),
	.Add2(\hps_0_h2f_axi_master_agent|Add2~0_combout ),
	.Add21(\hps_0_h2f_axi_master_agent|Add2~1_combout ),
	.Add22(\hps_0_h2f_axi_master_agent|Add2~2_combout ),
	.Add23(\hps_0_h2f_axi_master_agent|Add2~3_combout ),
	.write_cp_data_77(\hps_0_h2f_axi_master_agent|write_cp_data[77]~0_combout ),
	.write_cp_data_78(\hps_0_h2f_axi_master_agent|write_cp_data[78]~1_combout ),
	.write_cp_data_75(\hps_0_h2f_axi_master_agent|write_cp_data[75]~2_combout ),
	.write_cp_data_74(\hps_0_h2f_axi_master_agent|write_cp_data[74]~3_combout ),
	.write_cp_data_76(\hps_0_h2f_axi_master_agent|write_cp_data[76]~4_combout ),
	.WideNor0(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|WideNor0~0_combout ),
	.Equal14(\router|Equal14~1_combout ),
	.nxt_out_eop(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.src6_valid(\cmd_demux|src6_valid~1_combout ),
	.src_valid(\cmd_mux_006|src_valid~0_combout ),
	.cp_ready1(\wr_data_s1_agent|cp_ready~3_combout ),
	.in_data_reg_69(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.src_data_87(\cmd_mux_006|src_data[87]~combout ),
	.src_data_88(\cmd_mux_006|src_data[88]~combout ),
	.src_valid1(\cmd_mux_006|src_valid~1_combout ),
	.src_data_35(\cmd_mux_006|src_data[35]~combout ),
	.src_data_34(\cmd_mux_006|src_data[34]~combout ),
	.src_data_33(\cmd_mux_006|src_data[33]~combout ),
	.src_data_32(\cmd_mux_006|src_data[32]~combout ),
	.out_byte_cnt_reg_2(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_4(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_3(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_5(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_6(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.src_payload_0(\cmd_mux_006|src_payload[0]~combout ),
	.in_data_reg_105(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ),
	.in_data_reg_106(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ),
	.in_data_reg_107(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ),
	.in_data_reg_108(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ),
	.in_data_reg_109(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ),
	.in_data_reg_110(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ),
	.in_data_reg_111(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ),
	.in_data_reg_112(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ),
	.in_data_reg_113(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ),
	.in_data_reg_114(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ),
	.in_data_reg_115(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ),
	.in_data_reg_116(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ),
	.Selector3(\hps_0_h2f_axi_master_agent|Selector3~0_combout ),
	.Selector10(\hps_0_h2f_axi_master_agent|Selector10~1_combout ),
	.base_address_3(\hps_0_h2f_axi_master_agent|align_address_to_size|base_address[3]~0_combout ),
	.Selector4(\hps_0_h2f_axi_master_agent|Selector4~1_combout ),
	.Selector11(\hps_0_h2f_axi_master_agent|Selector11~1_combout ),
	.base_address_2(\hps_0_h2f_axi_master_agent|align_address_to_size|base_address[2]~1_combout ),
	.src_payload(\cmd_mux_006|src_payload~0_combout ),
	.src_data_82(\cmd_mux_006|src_data[82]~combout ),
	.src_data_81(\cmd_mux_006|src_data[81]~combout ),
	.src_data_105(\cmd_mux_006|src_data[105]~combout ),
	.src_data_106(\cmd_mux_006|src_data[106]~combout ),
	.src_data_107(\cmd_mux_006|src_data[107]~combout ),
	.src_data_108(\cmd_mux_006|src_data[108]~combout ),
	.src_data_109(\cmd_mux_006|src_data[109]~combout ),
	.src_data_110(\cmd_mux_006|src_data[110]~combout ),
	.src_data_111(\cmd_mux_006|src_data[111]~combout ),
	.src_data_112(\cmd_mux_006|src_data[112]~combout ),
	.src_data_113(\cmd_mux_006|src_data[113]~combout ),
	.src_data_114(\cmd_mux_006|src_data[114]~combout ),
	.src_data_115(\cmd_mux_006|src_data[115]~combout ),
	.src_data_116(\cmd_mux_006|src_data[116]~combout ),
	.src_data_86(\cmd_mux_006|src_data[86]~combout ),
	.Selector5(\hps_0_h2f_axi_master_agent|Selector5~1_combout ),
	.Selector12(\hps_0_h2f_axi_master_agent|Selector12~0_combout ),
	.out_data_1(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[1]~5_combout ),
	.src_data_80(\cmd_mux_006|src_data[80]~combout ),
	.out_data_0(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[0]~6_combout ),
	.Selector6(\hps_0_h2f_axi_master_agent|Selector6~0_combout ),
	.Selector13(\hps_0_h2f_axi_master_agent|Selector13~1_combout ),
	.src_data_79(\cmd_mux_006|src_data[79]~combout ),
	.clk_clk(clk_clk));

spw_babasu_altera_merlin_burst_adapter_2 data_i_s1_burst_adapter(
	.h2f_ARADDR_0(h2f_ARADDR_0),
	.h2f_ARADDR_1(h2f_ARADDR_1),
	.h2f_ARADDR_2(h2f_ARADDR_2),
	.h2f_ARADDR_3(h2f_ARADDR_3),
	.h2f_ARLEN_0(h2f_ARLEN_0),
	.nxt_in_ready(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.in_ready_hold(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.stateST_COMP_TRANS(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.out_valid_reg(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.in_narrow_reg(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.in_byteen_reg_3(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ),
	.in_byteen_reg_2(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ),
	.in_byteen_reg_1(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ),
	.in_byteen_reg_0(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ),
	.in_data_reg_68(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ),
	.cp_ready(\data_i_s1_agent|cp_ready~0_combout ),
	.stateST_UNCOMP_WR_SUBBURST(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.nxt_in_ready1(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.saved_grant_1(\cmd_mux_005|saved_grant[1]~q ),
	.Equal5(\router|Equal5~0_combout ),
	.saved_grant_0(\cmd_mux_005|saved_grant[0]~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.in_data_reg_0(in_data_reg_01),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_31),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_21),
	.in_data_reg_1(in_data_reg_1),
	.in_data_reg_2(in_data_reg_2),
	.in_data_reg_3(in_data_reg_3),
	.in_data_reg_4(in_data_reg_4),
	.in_data_reg_5(in_data_reg_5),
	.in_data_reg_6(in_data_reg_6),
	.in_data_reg_7(in_data_reg_7),
	.in_data_reg_8(in_data_reg_8),
	.Add2(\hps_0_h2f_axi_master_agent|Add2~0_combout ),
	.Add21(\hps_0_h2f_axi_master_agent|Add2~1_combout ),
	.Add22(\hps_0_h2f_axi_master_agent|Add2~2_combout ),
	.Add23(\hps_0_h2f_axi_master_agent|Add2~3_combout ),
	.Equal51(\router|Equal5~1_combout ),
	.write_cp_data_77(\hps_0_h2f_axi_master_agent|write_cp_data[77]~0_combout ),
	.write_cp_data_78(\hps_0_h2f_axi_master_agent|write_cp_data[78]~1_combout ),
	.write_cp_data_75(\hps_0_h2f_axi_master_agent|write_cp_data[75]~2_combout ),
	.write_cp_data_74(\hps_0_h2f_axi_master_agent|write_cp_data[74]~3_combout ),
	.write_cp_data_76(\hps_0_h2f_axi_master_agent|write_cp_data[76]~4_combout ),
	.WideNor0(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|WideNor0~0_combout ),
	.nxt_out_eop(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.src5_valid(\cmd_demux|src5_valid~1_combout ),
	.src_valid(\cmd_mux_005|src_valid~1_combout ),
	.cp_ready1(\data_i_s1_agent|cp_ready~3_combout ),
	.in_data_reg_69(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.src_data_87(\cmd_mux_005|src_data[87]~combout ),
	.src_data_88(\cmd_mux_005|src_data[88]~combout ),
	.src_valid1(\cmd_mux_005|src_valid~2_combout ),
	.src_data_35(\cmd_mux_005|src_data[35]~combout ),
	.src_data_34(\cmd_mux_005|src_data[34]~combout ),
	.src_data_33(\cmd_mux_005|src_data[33]~combout ),
	.src_data_32(\cmd_mux_005|src_data[32]~combout ),
	.out_byte_cnt_reg_2(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_3(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_4(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_5(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_6(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.src_payload_0(\cmd_mux_005|src_payload[0]~combout ),
	.in_data_reg_105(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ),
	.in_data_reg_106(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ),
	.in_data_reg_107(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ),
	.in_data_reg_108(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ),
	.in_data_reg_109(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ),
	.in_data_reg_110(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ),
	.in_data_reg_111(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ),
	.in_data_reg_112(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ),
	.in_data_reg_113(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ),
	.in_data_reg_114(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ),
	.in_data_reg_115(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ),
	.in_data_reg_116(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ),
	.Selector3(\hps_0_h2f_axi_master_agent|Selector3~0_combout ),
	.Selector10(\hps_0_h2f_axi_master_agent|Selector10~1_combout ),
	.base_address_3(\hps_0_h2f_axi_master_agent|align_address_to_size|base_address[3]~0_combout ),
	.Selector4(\hps_0_h2f_axi_master_agent|Selector4~1_combout ),
	.Selector11(\hps_0_h2f_axi_master_agent|Selector11~1_combout ),
	.base_address_2(\hps_0_h2f_axi_master_agent|align_address_to_size|base_address[2]~1_combout ),
	.src_payload(\cmd_mux_005|src_payload~0_combout ),
	.src_data_82(\cmd_mux_005|src_data[82]~combout ),
	.src_data_81(\cmd_mux_005|src_data[81]~combout ),
	.src_payload1(\cmd_mux_005|src_payload~1_combout ),
	.src_payload2(\cmd_mux_005|src_payload~2_combout ),
	.src_payload3(\cmd_mux_005|src_payload~3_combout ),
	.src_payload4(\cmd_mux_005|src_payload~4_combout ),
	.src_payload5(\cmd_mux_005|src_payload~5_combout ),
	.src_payload6(\cmd_mux_005|src_payload~6_combout ),
	.src_payload7(\cmd_mux_005|src_payload~7_combout ),
	.src_payload8(\cmd_mux_005|src_payload~8_combout ),
	.src_data_105(\cmd_mux_005|src_data[105]~combout ),
	.src_data_106(\cmd_mux_005|src_data[106]~combout ),
	.src_data_107(\cmd_mux_005|src_data[107]~combout ),
	.src_data_108(\cmd_mux_005|src_data[108]~combout ),
	.src_data_109(\cmd_mux_005|src_data[109]~combout ),
	.src_data_110(\cmd_mux_005|src_data[110]~combout ),
	.src_data_111(\cmd_mux_005|src_data[111]~combout ),
	.src_data_112(\cmd_mux_005|src_data[112]~combout ),
	.src_data_113(\cmd_mux_005|src_data[113]~combout ),
	.src_data_114(\cmd_mux_005|src_data[114]~combout ),
	.src_data_115(\cmd_mux_005|src_data[115]~combout ),
	.src_data_116(\cmd_mux_005|src_data[116]~combout ),
	.src_data_86(\cmd_mux_005|src_data[86]~combout ),
	.Selector5(\hps_0_h2f_axi_master_agent|Selector5~1_combout ),
	.Selector12(\hps_0_h2f_axi_master_agent|Selector12~0_combout ),
	.out_data_1(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[1]~5_combout ),
	.src_data_80(\cmd_mux_005|src_data[80]~combout ),
	.out_data_0(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[0]~6_combout ),
	.Selector6(\hps_0_h2f_axi_master_agent|Selector6~0_combout ),
	.Selector13(\hps_0_h2f_axi_master_agent|Selector13~1_combout ),
	.src_data_79(\cmd_mux_005|src_data[79]~combout ),
	.clk_clk(clk_clk));

spw_babasu_altera_merlin_burst_adapter_4 flags_s1_burst_adapter(
	.h2f_ARADDR_0(h2f_ARADDR_0),
	.h2f_ARADDR_1(h2f_ARADDR_1),
	.h2f_ARADDR_2(h2f_ARADDR_2),
	.h2f_ARADDR_3(h2f_ARADDR_3),
	.h2f_ARBURST_0(h2f_ARBURST_0),
	.h2f_ARBURST_1(h2f_ARBURST_1),
	.h2f_ARID_0(h2f_ARID_0),
	.h2f_ARID_1(h2f_ARID_1),
	.h2f_ARID_2(h2f_ARID_2),
	.h2f_ARID_3(h2f_ARID_3),
	.h2f_ARID_4(h2f_ARID_4),
	.h2f_ARID_5(h2f_ARID_5),
	.h2f_ARID_6(h2f_ARID_6),
	.h2f_ARID_7(h2f_ARID_7),
	.h2f_ARID_8(h2f_ARID_8),
	.h2f_ARID_9(h2f_ARID_9),
	.h2f_ARID_10(h2f_ARID_10),
	.h2f_ARID_11(h2f_ARID_11),
	.h2f_ARLEN_0(h2f_ARLEN_0),
	.Add5(\hps_0_h2f_axi_master_agent|Add5~1_sumout ),
	.Add51(\hps_0_h2f_axi_master_agent|Add5~5_sumout ),
	.in_ready_hold(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.in_data_reg_69(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.stateST_COMP_TRANS(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.mem_used_1(\flags_s1_agent_rsp_fifo|mem_used[1]~q ),
	.in_narrow_reg(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.cp_ready(\flags_s1_agent|cp_ready~0_combout ),
	.nxt_in_ready(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.out_valid_reg(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.stateST_UNCOMP_WR_SUBBURST(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.nxt_in_ready1(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.saved_grant_1(\cmd_mux_004|saved_grant[1]~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.Decoder1(\hps_0_h2f_axi_master_agent|Decoder1~0_combout ),
	.Add2(\hps_0_h2f_axi_master_agent|Add2~0_combout ),
	.Add21(\hps_0_h2f_axi_master_agent|Add2~1_combout ),
	.Add22(\hps_0_h2f_axi_master_agent|Add2~2_combout ),
	.Add23(\hps_0_h2f_axi_master_agent|Add2~3_combout ),
	.nxt_in_ready2(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ),
	.src_valid(\cmd_mux_004|src_valid~0_combout ),
	.nxt_out_eop(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.out_byte_cnt_reg_2(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.cp_ready1(\flags_s1_agent|cp_ready~1_combout ),
	.out_uncomp_byte_cnt_reg_6(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.out_uncomp_byte_cnt_reg_5(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_4(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_3(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.in_data_reg_105(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ),
	.in_data_reg_106(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ),
	.in_data_reg_107(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ),
	.in_data_reg_108(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ),
	.in_data_reg_109(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ),
	.in_data_reg_110(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ),
	.in_data_reg_111(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ),
	.in_data_reg_112(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ),
	.in_data_reg_113(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ),
	.in_data_reg_114(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ),
	.in_data_reg_115(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ),
	.in_data_reg_116(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ),
	.Selector10(\hps_0_h2f_axi_master_agent|Selector10~0_combout ),
	.Selector101(\hps_0_h2f_axi_master_agent|Selector10~1_combout ),
	.Selector11(\hps_0_h2f_axi_master_agent|Selector11~1_combout ),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_313),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_213),
	.Selector12(\hps_0_h2f_axi_master_agent|Selector12~0_combout ),
	.src_payload(\cmd_mux_004|src_payload~0_combout ),
	.src_payload1(\cmd_mux_004|src_payload~1_combout ),
	.src_payload2(\cmd_mux_004|src_payload~2_combout ),
	.Selector13(\hps_0_h2f_axi_master_agent|Selector13~1_combout ),
	.nxt_out_burstwrap_1(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_burstwrap[1]~0_combout ),
	.nxt_addr_2(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_addr[2]~2_combout ),
	.clk_clk(clk_clk));

spw_babasu_altera_merlin_burst_adapter_13 time_out_s1_burst_adapter(
	.h2f_ARADDR_0(h2f_ARADDR_0),
	.h2f_ARADDR_1(h2f_ARADDR_1),
	.h2f_ARADDR_2(h2f_ARADDR_2),
	.h2f_ARADDR_3(h2f_ARADDR_3),
	.h2f_ARBURST_0(h2f_ARBURST_0),
	.h2f_ARBURST_1(h2f_ARBURST_1),
	.h2f_ARID_0(h2f_ARID_0),
	.h2f_ARID_1(h2f_ARID_1),
	.h2f_ARID_2(h2f_ARID_2),
	.h2f_ARID_3(h2f_ARID_3),
	.h2f_ARID_4(h2f_ARID_4),
	.h2f_ARID_5(h2f_ARID_5),
	.h2f_ARID_6(h2f_ARID_6),
	.h2f_ARID_7(h2f_ARID_7),
	.h2f_ARID_8(h2f_ARID_8),
	.h2f_ARID_9(h2f_ARID_9),
	.h2f_ARID_10(h2f_ARID_10),
	.h2f_ARID_11(h2f_ARID_11),
	.h2f_ARLEN_0(h2f_ARLEN_0),
	.Add5(\hps_0_h2f_axi_master_agent|Add5~1_sumout ),
	.Add51(\hps_0_h2f_axi_master_agent|Add5~5_sumout ),
	.Add52(\hps_0_h2f_axi_master_agent|Add5~9_sumout ),
	.in_ready_hold(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.saved_grant_1(\cmd_mux_012|saved_grant[1]~q ),
	.stateST_COMP_TRANS(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.mem_used_1(\time_out_s1_agent_rsp_fifo|mem_used[1]~q ),
	.in_data_reg_69(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.in_narrow_reg(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.cp_ready(\time_out_s1_agent|cp_ready~0_combout ),
	.cp_ready1(\time_out_s1_agent|cp_ready~1_combout ),
	.nxt_out_eop(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.out_valid_reg(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.stateST_UNCOMP_WR_SUBBURST(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.nxt_in_ready(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.Decoder1(\hps_0_h2f_axi_master_agent|Decoder1~0_combout ),
	.Add2(\hps_0_h2f_axi_master_agent|Add2~0_combout ),
	.Add21(\hps_0_h2f_axi_master_agent|Add2~1_combout ),
	.Add22(\hps_0_h2f_axi_master_agent|Add2~2_combout ),
	.Add23(\hps_0_h2f_axi_master_agent|Add2~3_combout ),
	.nxt_in_ready1(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.src_valid(\cmd_mux_012|src_valid~0_combout ),
	.out_byte_cnt_reg_2(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.cp_ready2(\time_out_s1_agent|cp_ready~2_combout ),
	.out_uncomp_byte_cnt_reg_6(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.out_uncomp_byte_cnt_reg_5(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_4(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_3(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.in_data_reg_105(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ),
	.in_data_reg_106(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ),
	.in_data_reg_107(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ),
	.in_data_reg_108(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ),
	.in_data_reg_109(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ),
	.in_data_reg_110(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ),
	.in_data_reg_111(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ),
	.in_data_reg_112(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ),
	.in_data_reg_113(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ),
	.in_data_reg_114(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ),
	.in_data_reg_115(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ),
	.in_data_reg_116(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ),
	.Selector10(\hps_0_h2f_axi_master_agent|Selector10~0_combout ),
	.Selector101(\hps_0_h2f_axi_master_agent|Selector10~1_combout ),
	.Add3(\hps_0_h2f_axi_master_agent|Add3~1_combout ),
	.Add31(\hps_0_h2f_axi_master_agent|Add3~2_combout ),
	.Selector11(\hps_0_h2f_axi_master_agent|Selector11~0_combout ),
	.Selector111(\hps_0_h2f_axi_master_agent|Selector11~1_combout ),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_314),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_214),
	.Add32(\hps_0_h2f_axi_master_agent|Add3~3_combout ),
	.Selector12(\hps_0_h2f_axi_master_agent|Selector12~0_combout ),
	.src_payload(\cmd_mux_012|src_payload~0_combout ),
	.src_payload1(\cmd_mux_012|src_payload~1_combout ),
	.src_payload2(\cmd_mux_012|src_payload~2_combout ),
	.Selector13(\hps_0_h2f_axi_master_agent|Selector13~1_combout ),
	.nxt_out_burstwrap_1(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_burstwrap[1]~0_combout ),
	.nxt_addr_2(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_addr[2]~2_combout ),
	.clk_clk(clk_clk));

spw_babasu_altera_merlin_burst_adapter_11 tick_out_s1_burst_adapter(
	.h2f_ARADDR_0(h2f_ARADDR_0),
	.h2f_ARADDR_1(h2f_ARADDR_1),
	.h2f_ARADDR_2(h2f_ARADDR_2),
	.h2f_ARADDR_3(h2f_ARADDR_3),
	.h2f_ARBURST_0(h2f_ARBURST_0),
	.h2f_ARBURST_1(h2f_ARBURST_1),
	.h2f_ARID_0(h2f_ARID_0),
	.h2f_ARID_1(h2f_ARID_1),
	.h2f_ARID_2(h2f_ARID_2),
	.h2f_ARID_3(h2f_ARID_3),
	.h2f_ARID_4(h2f_ARID_4),
	.h2f_ARID_5(h2f_ARID_5),
	.h2f_ARID_6(h2f_ARID_6),
	.h2f_ARID_7(h2f_ARID_7),
	.h2f_ARID_8(h2f_ARID_8),
	.h2f_ARID_9(h2f_ARID_9),
	.h2f_ARID_10(h2f_ARID_10),
	.h2f_ARID_11(h2f_ARID_11),
	.h2f_ARLEN_0(h2f_ARLEN_0),
	.Add5(\hps_0_h2f_axi_master_agent|Add5~1_sumout ),
	.Add51(\hps_0_h2f_axi_master_agent|Add5~5_sumout ),
	.in_ready_hold(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.saved_grant_1(\cmd_mux_011|saved_grant[1]~q ),
	.stateST_COMP_TRANS(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.mem_used_1(\tick_out_s1_agent_rsp_fifo|mem_used[1]~q ),
	.in_data_reg_69(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.in_narrow_reg(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.cp_ready(\tick_out_s1_agent|cp_ready~0_combout ),
	.cp_ready1(\tick_out_s1_agent|cp_ready~1_combout ),
	.nxt_out_eop(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.out_valid_reg(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.stateST_UNCOMP_WR_SUBBURST(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.nxt_in_ready(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.Decoder1(\hps_0_h2f_axi_master_agent|Decoder1~0_combout ),
	.Add2(\hps_0_h2f_axi_master_agent|Add2~0_combout ),
	.Add21(\hps_0_h2f_axi_master_agent|Add2~1_combout ),
	.Add22(\hps_0_h2f_axi_master_agent|Add2~2_combout ),
	.Add23(\hps_0_h2f_axi_master_agent|Add2~3_combout ),
	.nxt_in_ready1(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.src_valid(\cmd_mux_011|src_valid~0_combout ),
	.out_byte_cnt_reg_2(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.cp_ready2(\tick_out_s1_agent|cp_ready~2_combout ),
	.out_uncomp_byte_cnt_reg_3(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_4(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_5(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_6(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.in_data_reg_105(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ),
	.in_data_reg_106(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ),
	.in_data_reg_107(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ),
	.in_data_reg_108(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ),
	.in_data_reg_109(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ),
	.in_data_reg_110(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ),
	.in_data_reg_111(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ),
	.in_data_reg_112(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ),
	.in_data_reg_113(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ),
	.in_data_reg_114(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ),
	.in_data_reg_115(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ),
	.in_data_reg_116(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ),
	.Selector10(\hps_0_h2f_axi_master_agent|Selector10~0_combout ),
	.Selector101(\hps_0_h2f_axi_master_agent|Selector10~1_combout ),
	.Selector11(\hps_0_h2f_axi_master_agent|Selector11~1_combout ),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_315),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_215),
	.Selector12(\hps_0_h2f_axi_master_agent|Selector12~0_combout ),
	.src_payload(\cmd_mux_011|src_payload~0_combout ),
	.src_payload1(\cmd_mux_011|src_payload~1_combout ),
	.src_payload2(\cmd_mux_011|src_payload~2_combout ),
	.Selector13(\hps_0_h2f_axi_master_agent|Selector13~1_combout ),
	.nxt_out_burstwrap_1(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_burstwrap[1]~0_combout ),
	.nxt_addr_2(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_addr[2]~2_combout ),
	.clk_clk(clk_clk));

spw_babasu_altera_merlin_burst_adapter_8 rx_empty_s1_burst_adapter(
	.h2f_ARADDR_0(h2f_ARADDR_0),
	.h2f_ARADDR_1(h2f_ARADDR_1),
	.h2f_ARADDR_2(h2f_ARADDR_2),
	.h2f_ARADDR_3(h2f_ARADDR_3),
	.h2f_ARBURST_0(h2f_ARBURST_0),
	.h2f_ARBURST_1(h2f_ARBURST_1),
	.h2f_ARID_0(h2f_ARID_0),
	.h2f_ARID_1(h2f_ARID_1),
	.h2f_ARID_2(h2f_ARID_2),
	.h2f_ARID_3(h2f_ARID_3),
	.h2f_ARID_4(h2f_ARID_4),
	.h2f_ARID_5(h2f_ARID_5),
	.h2f_ARID_6(h2f_ARID_6),
	.h2f_ARID_7(h2f_ARID_7),
	.h2f_ARID_8(h2f_ARID_8),
	.h2f_ARID_9(h2f_ARID_9),
	.h2f_ARID_10(h2f_ARID_10),
	.h2f_ARID_11(h2f_ARID_11),
	.h2f_ARLEN_0(h2f_ARLEN_0),
	.Add5(\hps_0_h2f_axi_master_agent|Add5~1_sumout ),
	.Add51(\hps_0_h2f_axi_master_agent|Add5~5_sumout ),
	.in_ready_hold(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.saved_grant_1(\cmd_mux_010|saved_grant[1]~q ),
	.stateST_COMP_TRANS(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.mem_used_1(\rx_empty_s1_agent_rsp_fifo|mem_used[1]~q ),
	.in_data_reg_69(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.in_narrow_reg(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.cp_ready(\rx_empty_s1_agent|cp_ready~0_combout ),
	.cp_ready1(\rx_empty_s1_agent|cp_ready~1_combout ),
	.nxt_out_eop(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.out_valid_reg(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.stateST_UNCOMP_WR_SUBBURST(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.nxt_in_ready(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.Decoder1(\hps_0_h2f_axi_master_agent|Decoder1~0_combout ),
	.Add2(\hps_0_h2f_axi_master_agent|Add2~0_combout ),
	.Add21(\hps_0_h2f_axi_master_agent|Add2~1_combout ),
	.Add22(\hps_0_h2f_axi_master_agent|Add2~2_combout ),
	.Add23(\hps_0_h2f_axi_master_agent|Add2~3_combout ),
	.src_valid(\cmd_mux_010|src_valid~0_combout ),
	.nxt_in_ready1(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.out_byte_cnt_reg_2(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.cp_ready2(\rx_empty_s1_agent|cp_ready~2_combout ),
	.out_uncomp_byte_cnt_reg_5(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_4(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_3(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_6(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.in_data_reg_105(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ),
	.in_data_reg_106(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ),
	.in_data_reg_107(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ),
	.in_data_reg_108(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ),
	.in_data_reg_109(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ),
	.in_data_reg_110(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ),
	.in_data_reg_111(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ),
	.in_data_reg_112(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ),
	.in_data_reg_113(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ),
	.in_data_reg_114(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ),
	.in_data_reg_115(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ),
	.in_data_reg_116(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ),
	.Selector10(\hps_0_h2f_axi_master_agent|Selector10~0_combout ),
	.Selector101(\hps_0_h2f_axi_master_agent|Selector10~1_combout ),
	.Selector11(\hps_0_h2f_axi_master_agent|Selector11~1_combout ),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_316),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_216),
	.Selector12(\hps_0_h2f_axi_master_agent|Selector12~0_combout ),
	.src_payload(\cmd_mux_010|src_payload~0_combout ),
	.src_payload1(\cmd_mux_010|src_payload~1_combout ),
	.src_payload2(\cmd_mux_010|src_payload~2_combout ),
	.Selector13(\hps_0_h2f_axi_master_agent|Selector13~1_combout ),
	.nxt_out_burstwrap_1(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_burstwrap[1]~0_combout ),
	.nxt_addr_2(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_addr[2]~2_combout ),
	.clk_clk(clk_clk));

spw_babasu_altera_merlin_burst_adapter_7 rd_data_s1_burst_adapter(
	.h2f_ARADDR_0(h2f_ARADDR_0),
	.h2f_ARADDR_1(h2f_ARADDR_1),
	.h2f_ARADDR_2(h2f_ARADDR_2),
	.h2f_ARADDR_3(h2f_ARADDR_3),
	.h2f_ARLEN_0(h2f_ARLEN_0),
	.nxt_in_ready(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.in_ready_hold(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.stateST_COMP_TRANS(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.out_valid_reg(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.in_narrow_reg(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.in_byteen_reg_3(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ),
	.in_byteen_reg_2(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ),
	.in_byteen_reg_1(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ),
	.in_byteen_reg_0(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ),
	.in_data_reg_68(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ),
	.cp_ready(\rd_data_s1_agent|cp_ready~0_combout ),
	.stateST_UNCOMP_WR_SUBBURST(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.nxt_in_ready1(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.saved_grant_1(\cmd_mux_009|saved_grant[1]~q ),
	.Equal9(\router|Equal9~0_combout ),
	.saved_grant_0(\cmd_mux_009|saved_grant[0]~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.in_data_reg_0(in_data_reg_04),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_34),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_24),
	.Add2(\hps_0_h2f_axi_master_agent|Add2~0_combout ),
	.Add21(\hps_0_h2f_axi_master_agent|Add2~1_combout ),
	.Add22(\hps_0_h2f_axi_master_agent|Add2~2_combout ),
	.Add23(\hps_0_h2f_axi_master_agent|Add2~3_combout ),
	.Equal5(\router|Equal5~1_combout ),
	.write_cp_data_77(\hps_0_h2f_axi_master_agent|write_cp_data[77]~0_combout ),
	.write_cp_data_78(\hps_0_h2f_axi_master_agent|write_cp_data[78]~1_combout ),
	.write_cp_data_75(\hps_0_h2f_axi_master_agent|write_cp_data[75]~2_combout ),
	.write_cp_data_74(\hps_0_h2f_axi_master_agent|write_cp_data[74]~3_combout ),
	.write_cp_data_76(\hps_0_h2f_axi_master_agent|write_cp_data[76]~4_combout ),
	.WideNor0(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|WideNor0~0_combout ),
	.nxt_out_eop(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.src9_valid(\cmd_demux|src9_valid~1_combout ),
	.src_valid(\cmd_mux_009|src_valid~0_combout ),
	.cp_ready1(\rd_data_s1_agent|cp_ready~3_combout ),
	.in_data_reg_69(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.src_data_87(\cmd_mux_009|src_data[87]~combout ),
	.src_data_88(\cmd_mux_009|src_data[88]~combout ),
	.src_valid1(\cmd_mux_009|src_valid~1_combout ),
	.src_data_35(\cmd_mux_009|src_data[35]~combout ),
	.src_data_34(\cmd_mux_009|src_data[34]~combout ),
	.src_data_33(\cmd_mux_009|src_data[33]~combout ),
	.src_data_32(\cmd_mux_009|src_data[32]~combout ),
	.out_byte_cnt_reg_2(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_4(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_3(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_5(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_6(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.src_payload_0(\cmd_mux_009|src_payload[0]~combout ),
	.in_data_reg_105(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ),
	.in_data_reg_106(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ),
	.in_data_reg_107(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ),
	.in_data_reg_108(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ),
	.in_data_reg_109(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ),
	.in_data_reg_110(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ),
	.in_data_reg_111(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ),
	.in_data_reg_112(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ),
	.in_data_reg_113(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ),
	.in_data_reg_114(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ),
	.in_data_reg_115(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ),
	.in_data_reg_116(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ),
	.Selector3(\hps_0_h2f_axi_master_agent|Selector3~0_combout ),
	.Selector10(\hps_0_h2f_axi_master_agent|Selector10~1_combout ),
	.base_address_3(\hps_0_h2f_axi_master_agent|align_address_to_size|base_address[3]~0_combout ),
	.Selector4(\hps_0_h2f_axi_master_agent|Selector4~1_combout ),
	.Selector11(\hps_0_h2f_axi_master_agent|Selector11~1_combout ),
	.base_address_2(\hps_0_h2f_axi_master_agent|align_address_to_size|base_address[2]~1_combout ),
	.src_payload(\cmd_mux_009|src_payload~0_combout ),
	.src_data_82(\cmd_mux_009|src_data[82]~combout ),
	.src_data_81(\cmd_mux_009|src_data[81]~combout ),
	.src_data_105(\cmd_mux_009|src_data[105]~combout ),
	.src_data_106(\cmd_mux_009|src_data[106]~combout ),
	.src_data_107(\cmd_mux_009|src_data[107]~combout ),
	.src_data_108(\cmd_mux_009|src_data[108]~combout ),
	.src_data_109(\cmd_mux_009|src_data[109]~combout ),
	.src_data_110(\cmd_mux_009|src_data[110]~combout ),
	.src_data_111(\cmd_mux_009|src_data[111]~combout ),
	.src_data_112(\cmd_mux_009|src_data[112]~combout ),
	.src_data_113(\cmd_mux_009|src_data[113]~combout ),
	.src_data_114(\cmd_mux_009|src_data[114]~combout ),
	.src_data_115(\cmd_mux_009|src_data[115]~combout ),
	.src_data_116(\cmd_mux_009|src_data[116]~combout ),
	.src_data_86(\cmd_mux_009|src_data[86]~combout ),
	.Selector5(\hps_0_h2f_axi_master_agent|Selector5~1_combout ),
	.Selector12(\hps_0_h2f_axi_master_agent|Selector12~0_combout ),
	.out_data_1(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[1]~5_combout ),
	.src_data_80(\cmd_mux_009|src_data[80]~combout ),
	.out_data_0(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[0]~6_combout ),
	.Selector6(\hps_0_h2f_axi_master_agent|Selector6~0_combout ),
	.Selector13(\hps_0_h2f_axi_master_agent|Selector13~1_combout ),
	.src_data_79(\cmd_mux_009|src_data[79]~combout ),
	.clk_clk(clk_clk));

spw_babasu_spw_babasu_mm_interconnect_0_cmd_mux cmd_mux(
	.h2f_WLAST_0(h2f_WLAST_0),
	.h2f_ARID_0(h2f_ARID_0),
	.h2f_ARID_1(h2f_ARID_1),
	.h2f_ARID_2(h2f_ARID_2),
	.h2f_ARID_3(h2f_ARID_3),
	.h2f_ARID_4(h2f_ARID_4),
	.h2f_ARID_5(h2f_ARID_5),
	.h2f_ARID_6(h2f_ARID_6),
	.h2f_ARID_7(h2f_ARID_7),
	.h2f_ARID_8(h2f_ARID_8),
	.h2f_ARID_9(h2f_ARID_9),
	.h2f_ARID_10(h2f_ARID_10),
	.h2f_ARID_11(h2f_ARID_11),
	.h2f_ARSIZE_0(h2f_ARSIZE_0),
	.h2f_ARSIZE_1(h2f_ARSIZE_1),
	.h2f_ARSIZE_2(h2f_ARSIZE_2),
	.h2f_AWID_0(h2f_AWID_0),
	.h2f_AWID_1(h2f_AWID_1),
	.h2f_AWID_2(h2f_AWID_2),
	.h2f_AWID_3(h2f_AWID_3),
	.h2f_AWID_4(h2f_AWID_4),
	.h2f_AWID_5(h2f_AWID_5),
	.h2f_AWID_6(h2f_AWID_6),
	.h2f_AWID_7(h2f_AWID_7),
	.h2f_AWID_8(h2f_AWID_8),
	.h2f_AWID_9(h2f_AWID_9),
	.h2f_AWID_10(h2f_AWID_10),
	.h2f_AWID_11(h2f_AWID_11),
	.h2f_AWSIZE_0(h2f_AWSIZE_0),
	.h2f_AWSIZE_1(h2f_AWSIZE_1),
	.h2f_AWSIZE_2(h2f_AWSIZE_2),
	.h2f_WDATA_0(h2f_WDATA_0),
	.h2f_WSTRB_0(h2f_WSTRB_0),
	.h2f_WSTRB_1(h2f_WSTRB_1),
	.h2f_WSTRB_2(h2f_WSTRB_2),
	.h2f_WSTRB_3(h2f_WSTRB_3),
	.nxt_in_ready(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~4_combout ),
	.saved_grant_1(\cmd_mux|saved_grant[1]~q ),
	.nxt_in_ready1(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.saved_grant_0(\cmd_mux|saved_grant[0]~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.src0_valid(\cmd_demux|src0_valid~1_combout ),
	.src0_valid1(\cmd_demux_001|src0_valid~0_combout ),
	.nxt_in_ready2(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ),
	.src_valid(\cmd_mux|src_valid~0_combout ),
	.src_payload_0(\cmd_mux|src_payload[0]~combout ),
	.src_data_87(\cmd_mux|src_data[87]~combout ),
	.src_data_88(\cmd_mux|src_data[88]~combout ),
	.src_data_35(\cmd_mux|src_data[35]~combout ),
	.src_data_34(\cmd_mux|src_data[34]~combout ),
	.src_data_33(\cmd_mux|src_data[33]~combout ),
	.src_data_32(\cmd_mux|src_data[32]~combout ),
	.Selector3(\hps_0_h2f_axi_master_agent|Selector3~0_combout ),
	.Selector10(\hps_0_h2f_axi_master_agent|Selector10~1_combout ),
	.Selector4(\hps_0_h2f_axi_master_agent|Selector4~1_combout ),
	.Selector11(\hps_0_h2f_axi_master_agent|Selector11~1_combout ),
	.src_payload(\cmd_mux|src_payload~0_combout ),
	.src_data_82(\cmd_mux|src_data[82]~combout ),
	.src_data_81(\cmd_mux|src_data[81]~combout ),
	.src_data_105(\cmd_mux|src_data[105]~combout ),
	.src_data_106(\cmd_mux|src_data[106]~combout ),
	.src_data_107(\cmd_mux|src_data[107]~combout ),
	.src_data_108(\cmd_mux|src_data[108]~combout ),
	.src_data_109(\cmd_mux|src_data[109]~combout ),
	.src_data_110(\cmd_mux|src_data[110]~combout ),
	.src_data_111(\cmd_mux|src_data[111]~combout ),
	.src_data_112(\cmd_mux|src_data[112]~combout ),
	.src_data_113(\cmd_mux|src_data[113]~combout ),
	.src_data_114(\cmd_mux|src_data[114]~combout ),
	.src_data_115(\cmd_mux|src_data[115]~combout ),
	.src_data_116(\cmd_mux|src_data[116]~combout ),
	.src_data_86(\cmd_mux|src_data[86]~combout ),
	.Selector5(\hps_0_h2f_axi_master_agent|Selector5~1_combout ),
	.Selector12(\hps_0_h2f_axi_master_agent|Selector12~0_combout ),
	.src_data_80(\cmd_mux|src_data[80]~combout ),
	.Selector6(\hps_0_h2f_axi_master_agent|Selector6~0_combout ),
	.Selector13(\hps_0_h2f_axi_master_agent|Selector13~1_combout ),
	.src_data_79(\cmd_mux|src_data[79]~combout ),
	.clk_clk(clk_clk));

spw_babasu_spw_babasu_mm_interconnect_0_cmd_demux_1 cmd_demux_001(
	.h2f_ARVALID_0(h2f_ARVALID_0),
	.h2f_ARADDR_4(h2f_ARADDR_4),
	.h2f_ARADDR_5(h2f_ARADDR_5),
	.h2f_ARADDR_6(h2f_ARADDR_6),
	.h2f_ARADDR_7(h2f_ARADDR_7),
	.h2f_ARADDR_8(h2f_ARADDR_8),
	.nxt_in_ready(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.nxt_in_ready1(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.nxt_in_ready2(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~4_combout ),
	.nxt_in_ready3(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.nxt_in_ready4(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.nxt_in_ready5(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.nxt_in_ready6(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.nxt_in_ready7(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ),
	.nxt_in_ready8(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.nxt_in_ready9(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.has_pending_responses(\hps_0_h2f_axi_master_rd_limiter|has_pending_responses~q ),
	.last_channel_6(\hps_0_h2f_axi_master_rd_limiter|last_channel[6]~q ),
	.Equal6(\router_001|Equal6~0_combout ),
	.saved_grant_1(\cmd_mux_008|saved_grant[1]~q ),
	.stateST_COMP_TRANS(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.cp_ready(\data_o_s1_agent|cp_ready~1_combout ),
	.nxt_out_eop(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.src_channel(\router_001|src_channel~0_combout ),
	.nxt_in_ready10(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.saved_grant_11(\cmd_mux_011|saved_grant[1]~q ),
	.stateST_COMP_TRANS1(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.cp_ready1(\tick_out_s1_agent|cp_ready~1_combout ),
	.nxt_out_eop1(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.last_cycle(\cmd_mux_011|last_cycle~0_combout ),
	.nxt_in_ready11(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.saved_grant_12(\cmd_mux_012|saved_grant[1]~q ),
	.stateST_COMP_TRANS2(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.cp_ready2(\time_out_s1_agent|cp_ready~1_combout ),
	.nxt_out_eop2(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.last_cycle1(\cmd_mux_012|last_cycle~0_combout ),
	.nxt_in_ready12(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.nxt_in_ready13(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.saved_grant_13(\cmd_mux_001|saved_grant[1]~q ),
	.src_channel_1(\router_001|src_channel[1]~1_combout ),
	.WideOr0(\cmd_demux_001|WideOr0~0_combout ),
	.nxt_in_ready14(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.saved_grant_14(\cmd_mux_015|saved_grant[1]~q ),
	.Equal15(\router_001|Equal15~0_combout ),
	.nxt_in_ready15(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.Equal16(\router_001|Equal16~0_combout ),
	.saved_grant_15(\cmd_mux_016|saved_grant[1]~q ),
	.WideOr01(\cmd_demux_001|WideOr0~1_combout ),
	.nxt_in_ready16(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.saved_grant_16(\cmd_mux_013|saved_grant[1]~q ),
	.src_channel_13(\router_001|src_channel[13]~2_combout ),
	.nxt_in_ready17(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.saved_grant_17(\cmd_mux_014|saved_grant[1]~q ),
	.Equal14(\router_001|Equal14~0_combout ),
	.WideOr02(\cmd_demux_001|WideOr0~2_combout ),
	.Equal3(\router_001|Equal3~0_combout ),
	.saved_grant_18(\cmd_mux_003|saved_grant[1]~q ),
	.stateST_COMP_TRANS3(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.cp_ready3(\currentstate_s1_agent|cp_ready~1_combout ),
	.nxt_out_eop3(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.nxt_in_ready18(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.nxt_in_ready19(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.saved_grant_19(\cmd_mux_005|saved_grant[1]~q ),
	.nxt_in_ready20(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.saved_grant_110(\cmd_mux_009|saved_grant[1]~q ),
	.saved_grant_111(\cmd_mux_010|saved_grant[1]~q ),
	.Equal10(\router_001|Equal10~0_combout ),
	.stateST_COMP_TRANS4(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.cp_ready4(\rx_empty_s1_agent|cp_ready~1_combout ),
	.nxt_out_eop4(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.nxt_in_ready21(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.saved_grant_112(\cmd_mux|saved_grant[1]~q ),
	.nxt_in_ready22(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.src_channel_0(\router_001|src_channel[0]~3_combout ),
	.nxt_in_ready23(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.nxt_in_ready24(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.nxt_in_ready25(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.saved_grant_113(\cmd_mux_004|saved_grant[1]~q ),
	.nxt_in_ready26(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.saved_grant_114(\cmd_mux_007|saved_grant[1]~q ),
	.nxt_in_ready27(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.saved_grant_115(\cmd_mux_002|saved_grant[1]~q ),
	.nxt_in_ready28(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.saved_grant_116(\cmd_mux_006|saved_grant[1]~q ),
	.WideOr03(\cmd_demux_001|WideOr0~6_combout ),
	.last_channel_1(\hps_0_h2f_axi_master_rd_limiter|last_channel[1]~q ),
	.src1_valid(\cmd_demux_001|src1_valid~0_combout ),
	.last_channel_15(\hps_0_h2f_axi_master_rd_limiter|last_channel[15]~q ),
	.src15_valid(\cmd_demux_001|src15_valid~0_combout ),
	.src15_valid1(\cmd_demux_001|src15_valid~1_combout ),
	.last_channel_16(\hps_0_h2f_axi_master_rd_limiter|last_channel[16]~q ),
	.src16_valid(\cmd_demux_001|src16_valid~0_combout ),
	.src16_valid1(\cmd_demux_001|src16_valid~1_combout ),
	.last_channel_14(\hps_0_h2f_axi_master_rd_limiter|last_channel[14]~q ),
	.src14_valid(\cmd_demux_001|src14_valid~0_combout ),
	.src14_valid1(\cmd_demux_001|src14_valid~1_combout ),
	.Equal9(\router_001|Equal9~0_combout ),
	.last_channel_9(\hps_0_h2f_axi_master_rd_limiter|last_channel[9]~q ),
	.src9_valid(\cmd_demux_001|src9_valid~0_combout ),
	.src9_valid1(\cmd_demux_001|src9_valid~1_combout ),
	.last_channel_0(\hps_0_h2f_axi_master_rd_limiter|last_channel[0]~q ),
	.src0_valid(\cmd_demux_001|src0_valid~0_combout ),
	.src_channel_2(\router_001|src_channel[2]~4_combout ),
	.last_channel_2(\hps_0_h2f_axi_master_rd_limiter|last_channel[2]~q ),
	.src2_valid(\cmd_demux_001|src2_valid~0_combout ),
	.src2_valid1(\cmd_demux_001|src2_valid~1_combout ),
	.src6_valid(\cmd_demux_001|src6_valid~0_combout ),
	.src6_valid1(\cmd_demux_001|src6_valid~1_combout ));

spw_babasu_spw_babasu_mm_interconnect_0_cmd_demux cmd_demux(
	.h2f_AWVALID_0(h2f_AWVALID_0),
	.h2f_WVALID_0(h2f_WVALID_0),
	.nxt_in_ready(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.nxt_in_ready1(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.nxt_in_ready2(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~4_combout ),
	.nxt_in_ready3(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.nxt_in_ready4(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.nxt_in_ready5(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.nxt_in_ready6(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.nxt_in_ready7(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ),
	.nxt_in_ready8(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.nxt_in_ready9(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.nxt_in_ready10(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.nxt_in_ready11(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.nxt_in_ready12(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.nxt_in_ready13(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.nxt_in_ready14(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.nxt_in_ready15(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.nxt_in_ready16(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.nxt_in_ready17(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.nxt_in_ready18(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.nxt_in_ready19(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.write_addr_data_both_valid(\hps_0_h2f_axi_master_agent|write_addr_data_both_valid~combout ),
	.has_pending_responses(\hps_0_h2f_axi_master_wr_limiter|has_pending_responses~q ),
	.out_data_8(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[8]~0_combout ),
	.out_data_5(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[5]~1_combout ),
	.out_data_4(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[4]~2_combout ),
	.out_data_7(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[7]~3_combout ),
	.out_data_6(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[6]~4_combout ),
	.Equal5(\router|Equal5~0_combout ),
	.Equal14(\router|Equal14~0_combout ),
	.last_channel_6(\hps_0_h2f_axi_master_wr_limiter|last_channel[6]~q ),
	.Equal16(\router|Equal16~0_combout ),
	.Equal13(\router|Equal13~0_combout ),
	.Equal15(\router|Equal15~0_combout ),
	.saved_grant_0(\cmd_mux_015|saved_grant[0]~q ),
	.Equal161(\router|Equal16~1_combout ),
	.saved_grant_01(\cmd_mux_016|saved_grant[0]~q ),
	.WideOr0(\cmd_demux|WideOr0~0_combout ),
	.saved_grant_02(\cmd_mux_013|saved_grant[0]~q ),
	.saved_grant_03(\cmd_mux_014|saved_grant[0]~q ),
	.WideOr01(\cmd_demux|WideOr0~1_combout ),
	.saved_grant_04(\cmd_mux_006|saved_grant[0]~q ),
	.Equal9(\router|Equal9~0_combout ),
	.saved_grant_05(\cmd_mux_009|saved_grant[0]~q ),
	.WideOr02(\cmd_demux|WideOr0~2_combout ),
	.saved_grant_06(\cmd_mux|saved_grant[0]~q ),
	.saved_grant_07(\cmd_mux_001|saved_grant[0]~q ),
	.WideOr03(\cmd_demux|WideOr0~3_combout ),
	.saved_grant_08(\cmd_mux_002|saved_grant[0]~q ),
	.saved_grant_09(\cmd_mux_005|saved_grant[0]~q ),
	.WideOr04(\cmd_demux|WideOr0~4_combout ),
	.WideOr05(\cmd_demux|WideOr0~5_combout ),
	.last_channel_1(\hps_0_h2f_axi_master_wr_limiter|last_channel[1]~q ),
	.src1_valid(\cmd_demux|src1_valid~0_combout ),
	.src1_valid1(\cmd_demux|src1_valid~1_combout ),
	.src1_valid2(\cmd_demux|src1_valid~2_combout ),
	.last_channel_15(\hps_0_h2f_axi_master_wr_limiter|last_channel[15]~q ),
	.src15_valid(\cmd_demux|src15_valid~0_combout ),
	.src15_valid1(\cmd_demux|src15_valid~1_combout ),
	.src15_valid2(\cmd_demux|src15_valid~2_combout ),
	.last_channel_16(\hps_0_h2f_axi_master_wr_limiter|last_channel[16]~q ),
	.src16_valid(\cmd_demux|src16_valid~0_combout ),
	.src16_valid1(\cmd_demux|src16_valid~1_combout ),
	.src16_valid2(\cmd_demux|src16_valid~2_combout ),
	.last_channel_13(\hps_0_h2f_axi_master_wr_limiter|last_channel[13]~q ),
	.src13_valid(\cmd_demux|src13_valid~0_combout ),
	.src13_valid1(\cmd_demux|src13_valid~1_combout ),
	.src13_valid2(\cmd_demux|src13_valid~2_combout ),
	.last_channel_14(\hps_0_h2f_axi_master_wr_limiter|last_channel[14]~q ),
	.src14_valid(\cmd_demux|src14_valid~0_combout ),
	.src14_valid1(\cmd_demux|src14_valid~1_combout ),
	.src14_valid2(\cmd_demux|src14_valid~2_combout ),
	.last_channel_5(\hps_0_h2f_axi_master_wr_limiter|last_channel[5]~q ),
	.src5_valid(\cmd_demux|src5_valid~0_combout ),
	.src5_valid1(\cmd_demux|src5_valid~1_combout ),
	.src5_valid2(\cmd_demux|src5_valid~2_combout ),
	.last_channel_9(\hps_0_h2f_axi_master_wr_limiter|last_channel[9]~q ),
	.src9_valid(\cmd_demux|src9_valid~0_combout ),
	.src9_valid1(\cmd_demux|src9_valid~1_combout ),
	.src9_valid2(\cmd_demux|src9_valid~2_combout ),
	.last_channel_0(\hps_0_h2f_axi_master_wr_limiter|last_channel[0]~q ),
	.src0_valid(\cmd_demux|src0_valid~1_combout ),
	.last_channel_2(\hps_0_h2f_axi_master_wr_limiter|last_channel[2]~q ),
	.src2_valid(\cmd_demux|src2_valid~0_combout ),
	.src2_valid1(\cmd_demux|src2_valid~1_combout ),
	.src2_valid2(\cmd_demux|src2_valid~2_combout ),
	.src6_valid(\cmd_demux|src6_valid~0_combout ),
	.src6_valid1(\cmd_demux|src6_valid~1_combout ),
	.src6_valid2(\cmd_demux|src6_valid~2_combout ));

spw_babasu_altera_merlin_burst_adapter_9 spill_enable_s1_burst_adapter(
	.h2f_ARADDR_0(h2f_ARADDR_0),
	.h2f_ARADDR_1(h2f_ARADDR_1),
	.h2f_ARADDR_2(h2f_ARADDR_2),
	.h2f_ARADDR_3(h2f_ARADDR_3),
	.h2f_ARLEN_0(h2f_ARLEN_0),
	.nxt_in_ready(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ),
	.in_ready_hold(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.stateST_COMP_TRANS(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.out_valid_reg(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\spill_enable_s1_agent_rsp_fifo|mem_used[1]~q ),
	.in_narrow_reg(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.in_byteen_reg_3(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ),
	.in_byteen_reg_2(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ),
	.in_byteen_reg_1(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ),
	.in_byteen_reg_0(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ),
	.in_data_reg_68(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ),
	.cp_ready(\spill_enable_s1_agent|cp_ready~0_combout ),
	.stateST_UNCOMP_WR_SUBBURST(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.nxt_in_ready1(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.saved_grant_1(\cmd_mux_016|saved_grant[1]~q ),
	.saved_grant_0(\cmd_mux_016|saved_grant[0]~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.in_data_reg_0(in_data_reg_05),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_35),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_25),
	.Add2(\hps_0_h2f_axi_master_agent|Add2~0_combout ),
	.Add21(\hps_0_h2f_axi_master_agent|Add2~1_combout ),
	.Add22(\hps_0_h2f_axi_master_agent|Add2~2_combout ),
	.Add23(\hps_0_h2f_axi_master_agent|Add2~3_combout ),
	.write_cp_data_77(\hps_0_h2f_axi_master_agent|write_cp_data[77]~0_combout ),
	.write_cp_data_78(\hps_0_h2f_axi_master_agent|write_cp_data[78]~1_combout ),
	.write_cp_data_75(\hps_0_h2f_axi_master_agent|write_cp_data[75]~2_combout ),
	.write_cp_data_74(\hps_0_h2f_axi_master_agent|write_cp_data[74]~3_combout ),
	.write_cp_data_76(\hps_0_h2f_axi_master_agent|write_cp_data[76]~4_combout ),
	.WideNor0(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|WideNor0~0_combout ),
	.nxt_out_eop(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.src_valid(\cmd_mux_016|src_valid~0_combout ),
	.src_valid1(\cmd_mux_016|src_valid~1_combout ),
	.WideOr1(\cmd_mux_016|WideOr1~combout ),
	.cp_ready1(\spill_enable_s1_agent|cp_ready~1_combout ),
	.cp_ready2(\spill_enable_s1_agent|cp_ready~2_combout ),
	.in_data_reg_69(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.src_data_87(\cmd_mux_016|src_data[87]~combout ),
	.src_data_88(\cmd_mux_016|src_data[88]~combout ),
	.src_data_35(\cmd_mux_016|src_data[35]~combout ),
	.src_data_34(\cmd_mux_016|src_data[34]~combout ),
	.src_data_33(\cmd_mux_016|src_data[33]~combout ),
	.src_data_32(\cmd_mux_016|src_data[32]~combout ),
	.out_byte_cnt_reg_2(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_5(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_4(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_3(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_6(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.src_payload_0(\cmd_mux_016|src_payload[0]~combout ),
	.in_data_reg_105(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ),
	.in_data_reg_106(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ),
	.in_data_reg_107(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ),
	.in_data_reg_108(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ),
	.in_data_reg_109(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ),
	.in_data_reg_110(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ),
	.in_data_reg_111(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ),
	.in_data_reg_112(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ),
	.in_data_reg_113(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ),
	.in_data_reg_114(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ),
	.in_data_reg_115(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ),
	.in_data_reg_116(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ),
	.Selector3(\hps_0_h2f_axi_master_agent|Selector3~0_combout ),
	.Selector10(\hps_0_h2f_axi_master_agent|Selector10~1_combout ),
	.base_address_3(\hps_0_h2f_axi_master_agent|align_address_to_size|base_address[3]~0_combout ),
	.Selector4(\hps_0_h2f_axi_master_agent|Selector4~1_combout ),
	.Selector11(\hps_0_h2f_axi_master_agent|Selector11~1_combout ),
	.base_address_2(\hps_0_h2f_axi_master_agent|align_address_to_size|base_address[2]~1_combout ),
	.src_payload(\cmd_mux_016|src_payload~0_combout ),
	.src_data_82(\cmd_mux_016|src_data[82]~combout ),
	.src_data_81(\cmd_mux_016|src_data[81]~combout ),
	.src_data_105(\cmd_mux_016|src_data[105]~combout ),
	.src_data_106(\cmd_mux_016|src_data[106]~combout ),
	.src_data_107(\cmd_mux_016|src_data[107]~combout ),
	.src_data_108(\cmd_mux_016|src_data[108]~combout ),
	.src_data_109(\cmd_mux_016|src_data[109]~combout ),
	.src_data_110(\cmd_mux_016|src_data[110]~combout ),
	.src_data_111(\cmd_mux_016|src_data[111]~combout ),
	.src_data_112(\cmd_mux_016|src_data[112]~combout ),
	.src_data_113(\cmd_mux_016|src_data[113]~combout ),
	.src_data_114(\cmd_mux_016|src_data[114]~combout ),
	.src_data_115(\cmd_mux_016|src_data[115]~combout ),
	.src_data_116(\cmd_mux_016|src_data[116]~combout ),
	.src_data_86(\cmd_mux_016|src_data[86]~combout ),
	.Selector5(\hps_0_h2f_axi_master_agent|Selector5~1_combout ),
	.Selector12(\hps_0_h2f_axi_master_agent|Selector12~0_combout ),
	.out_data_1(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[1]~5_combout ),
	.src_data_80(\cmd_mux_016|src_data[80]~combout ),
	.out_data_0(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[0]~6_combout ),
	.Selector6(\hps_0_h2f_axi_master_agent|Selector6~0_combout ),
	.Selector13(\hps_0_h2f_axi_master_agent|Selector13~1_combout ),
	.src_data_79(\cmd_mux_016|src_data[79]~combout ),
	.clk_clk(clk_clk));

spw_babasu_altera_merlin_burst_adapter_14 tx_clk_div_s1_burst_adapter(
	.h2f_ARADDR_0(h2f_ARADDR_0),
	.h2f_ARADDR_1(h2f_ARADDR_1),
	.h2f_ARADDR_2(h2f_ARADDR_2),
	.h2f_ARADDR_3(h2f_ARADDR_3),
	.h2f_ARLEN_0(h2f_ARLEN_0),
	.nxt_in_ready(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.in_ready_hold(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.stateST_COMP_TRANS(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.out_valid_reg(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.in_narrow_reg(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.in_byteen_reg_3(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ),
	.in_byteen_reg_2(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ),
	.in_byteen_reg_1(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ),
	.in_byteen_reg_0(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ),
	.in_data_reg_68(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ),
	.cp_ready(\tx_clk_div_s1_agent|cp_ready~0_combout ),
	.stateST_UNCOMP_WR_SUBBURST(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.nxt_in_ready1(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.saved_grant_1(\cmd_mux_015|saved_grant[1]~q ),
	.Equal15(\router|Equal15~0_combout ),
	.saved_grant_0(\cmd_mux_015|saved_grant[0]~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.in_data_reg_0(in_data_reg_08),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_38),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_28),
	.in_data_reg_1(in_data_reg_12),
	.in_data_reg_2(in_data_reg_22),
	.in_data_reg_3(in_data_reg_32),
	.in_data_reg_4(in_data_reg_42),
	.in_data_reg_5(in_data_reg_52),
	.in_data_reg_6(in_data_reg_62),
	.Add2(\hps_0_h2f_axi_master_agent|Add2~0_combout ),
	.Add21(\hps_0_h2f_axi_master_agent|Add2~1_combout ),
	.Add22(\hps_0_h2f_axi_master_agent|Add2~2_combout ),
	.Add23(\hps_0_h2f_axi_master_agent|Add2~3_combout ),
	.write_cp_data_77(\hps_0_h2f_axi_master_agent|write_cp_data[77]~0_combout ),
	.write_cp_data_78(\hps_0_h2f_axi_master_agent|write_cp_data[78]~1_combout ),
	.write_cp_data_75(\hps_0_h2f_axi_master_agent|write_cp_data[75]~2_combout ),
	.write_cp_data_74(\hps_0_h2f_axi_master_agent|write_cp_data[74]~3_combout ),
	.write_cp_data_76(\hps_0_h2f_axi_master_agent|write_cp_data[76]~4_combout ),
	.WideNor0(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|WideNor0~0_combout ),
	.nxt_out_eop(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.Equal151(\router|Equal15~1_combout ),
	.src15_valid(\cmd_demux|src15_valid~1_combout ),
	.src_valid(\cmd_mux_015|src_valid~0_combout ),
	.cp_ready1(\tx_clk_div_s1_agent|cp_ready~3_combout ),
	.in_data_reg_69(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.src_data_87(\cmd_mux_015|src_data[87]~combout ),
	.src_data_88(\cmd_mux_015|src_data[88]~combout ),
	.src_valid1(\cmd_mux_015|src_valid~1_combout ),
	.src_data_35(\cmd_mux_015|src_data[35]~combout ),
	.src_data_34(\cmd_mux_015|src_data[34]~combout ),
	.src_data_33(\cmd_mux_015|src_data[33]~combout ),
	.src_data_32(\cmd_mux_015|src_data[32]~combout ),
	.out_byte_cnt_reg_2(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_4(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_3(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_5(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_6(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.src_payload_0(\cmd_mux_015|src_payload[0]~combout ),
	.in_data_reg_105(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ),
	.in_data_reg_106(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ),
	.in_data_reg_107(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ),
	.in_data_reg_108(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ),
	.in_data_reg_109(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ),
	.in_data_reg_110(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ),
	.in_data_reg_111(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ),
	.in_data_reg_112(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ),
	.in_data_reg_113(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ),
	.in_data_reg_114(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ),
	.in_data_reg_115(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ),
	.in_data_reg_116(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ),
	.Selector3(\hps_0_h2f_axi_master_agent|Selector3~0_combout ),
	.Selector10(\hps_0_h2f_axi_master_agent|Selector10~1_combout ),
	.base_address_3(\hps_0_h2f_axi_master_agent|align_address_to_size|base_address[3]~0_combout ),
	.Selector4(\hps_0_h2f_axi_master_agent|Selector4~1_combout ),
	.Selector11(\hps_0_h2f_axi_master_agent|Selector11~1_combout ),
	.base_address_2(\hps_0_h2f_axi_master_agent|align_address_to_size|base_address[2]~1_combout ),
	.src_payload(\cmd_mux_015|src_payload~0_combout ),
	.src_data_82(\cmd_mux_015|src_data[82]~combout ),
	.src_data_81(\cmd_mux_015|src_data[81]~combout ),
	.src_payload1(\cmd_mux_015|src_payload~1_combout ),
	.src_payload2(\cmd_mux_015|src_payload~2_combout ),
	.src_payload3(\cmd_mux_015|src_payload~3_combout ),
	.src_payload4(\cmd_mux_015|src_payload~4_combout ),
	.src_payload5(\cmd_mux_015|src_payload~5_combout ),
	.src_payload6(\cmd_mux_015|src_payload~6_combout ),
	.src_data_105(\cmd_mux_015|src_data[105]~combout ),
	.src_data_106(\cmd_mux_015|src_data[106]~combout ),
	.src_data_107(\cmd_mux_015|src_data[107]~combout ),
	.src_data_108(\cmd_mux_015|src_data[108]~combout ),
	.src_data_109(\cmd_mux_015|src_data[109]~combout ),
	.src_data_110(\cmd_mux_015|src_data[110]~combout ),
	.src_data_111(\cmd_mux_015|src_data[111]~combout ),
	.src_data_112(\cmd_mux_015|src_data[112]~combout ),
	.src_data_113(\cmd_mux_015|src_data[113]~combout ),
	.src_data_114(\cmd_mux_015|src_data[114]~combout ),
	.src_data_115(\cmd_mux_015|src_data[115]~combout ),
	.src_data_116(\cmd_mux_015|src_data[116]~combout ),
	.src_data_86(\cmd_mux_015|src_data[86]~combout ),
	.Selector5(\hps_0_h2f_axi_master_agent|Selector5~1_combout ),
	.Selector12(\hps_0_h2f_axi_master_agent|Selector12~0_combout ),
	.out_data_1(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[1]~5_combout ),
	.src_data_80(\cmd_mux_015|src_data[80]~combout ),
	.out_data_0(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[0]~6_combout ),
	.Selector6(\hps_0_h2f_axi_master_agent|Selector6~0_combout ),
	.Selector13(\hps_0_h2f_axi_master_agent|Selector13~1_combout ),
	.src_data_79(\cmd_mux_015|src_data[79]~combout ),
	.clk_clk(clk_clk));

spw_babasu_altera_merlin_burst_adapter_12 time_in_s1_burst_adapter(
	.h2f_ARADDR_0(h2f_ARADDR_0),
	.h2f_ARADDR_1(h2f_ARADDR_1),
	.h2f_ARADDR_2(h2f_ARADDR_2),
	.h2f_ARADDR_3(h2f_ARADDR_3),
	.h2f_ARLEN_0(h2f_ARLEN_0),
	.nxt_in_ready(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.in_ready_hold(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.stateST_COMP_TRANS(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.out_valid_reg(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.in_narrow_reg(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.in_byteen_reg_3(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ),
	.in_byteen_reg_2(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ),
	.in_byteen_reg_1(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ),
	.in_byteen_reg_0(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ),
	.in_data_reg_68(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ),
	.cp_ready(\time_in_s1_agent|cp_ready~0_combout ),
	.stateST_UNCOMP_WR_SUBBURST(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.nxt_in_ready1(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.saved_grant_1(\cmd_mux_014|saved_grant[1]~q ),
	.Equal13(\router|Equal13~0_combout ),
	.saved_grant_0(\cmd_mux_014|saved_grant[0]~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.in_data_reg_0(in_data_reg_07),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_37),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_27),
	.in_data_reg_1(in_data_reg_11),
	.in_data_reg_2(in_data_reg_21),
	.in_data_reg_3(in_data_reg_31),
	.in_data_reg_4(in_data_reg_41),
	.in_data_reg_5(in_data_reg_51),
	.in_data_reg_6(in_data_reg_61),
	.in_data_reg_7(in_data_reg_71),
	.Add2(\hps_0_h2f_axi_master_agent|Add2~0_combout ),
	.Add21(\hps_0_h2f_axi_master_agent|Add2~1_combout ),
	.Add22(\hps_0_h2f_axi_master_agent|Add2~2_combout ),
	.Add23(\hps_0_h2f_axi_master_agent|Add2~3_combout ),
	.write_cp_data_77(\hps_0_h2f_axi_master_agent|write_cp_data[77]~0_combout ),
	.write_cp_data_78(\hps_0_h2f_axi_master_agent|write_cp_data[78]~1_combout ),
	.write_cp_data_75(\hps_0_h2f_axi_master_agent|write_cp_data[75]~2_combout ),
	.write_cp_data_74(\hps_0_h2f_axi_master_agent|write_cp_data[74]~3_combout ),
	.write_cp_data_76(\hps_0_h2f_axi_master_agent|write_cp_data[76]~4_combout ),
	.WideNor0(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|WideNor0~0_combout ),
	.nxt_out_eop(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.Equal14(\router|Equal14~1_combout ),
	.src14_valid(\cmd_demux|src14_valid~1_combout ),
	.src_valid(\cmd_mux_014|src_valid~0_combout ),
	.cp_ready1(\time_in_s1_agent|cp_ready~3_combout ),
	.in_data_reg_69(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.src_data_87(\cmd_mux_014|src_data[87]~combout ),
	.src_data_88(\cmd_mux_014|src_data[88]~combout ),
	.src_valid1(\cmd_mux_014|src_valid~1_combout ),
	.src_data_35(\cmd_mux_014|src_data[35]~combout ),
	.src_data_34(\cmd_mux_014|src_data[34]~combout ),
	.src_data_33(\cmd_mux_014|src_data[33]~combout ),
	.src_data_32(\cmd_mux_014|src_data[32]~combout ),
	.out_byte_cnt_reg_2(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_5(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_4(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_3(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_6(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.src_payload_0(\cmd_mux_014|src_payload[0]~combout ),
	.in_data_reg_105(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ),
	.in_data_reg_106(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ),
	.in_data_reg_107(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ),
	.in_data_reg_108(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ),
	.in_data_reg_109(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ),
	.in_data_reg_110(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ),
	.in_data_reg_111(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ),
	.in_data_reg_112(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ),
	.in_data_reg_113(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ),
	.in_data_reg_114(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ),
	.in_data_reg_115(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ),
	.in_data_reg_116(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ),
	.Selector3(\hps_0_h2f_axi_master_agent|Selector3~0_combout ),
	.Selector10(\hps_0_h2f_axi_master_agent|Selector10~1_combout ),
	.base_address_3(\hps_0_h2f_axi_master_agent|align_address_to_size|base_address[3]~0_combout ),
	.Selector4(\hps_0_h2f_axi_master_agent|Selector4~1_combout ),
	.Selector11(\hps_0_h2f_axi_master_agent|Selector11~1_combout ),
	.base_address_2(\hps_0_h2f_axi_master_agent|align_address_to_size|base_address[2]~1_combout ),
	.src_payload(\cmd_mux_014|src_payload~0_combout ),
	.src_data_82(\cmd_mux_014|src_data[82]~combout ),
	.src_data_81(\cmd_mux_014|src_data[81]~combout ),
	.src_payload1(\cmd_mux_014|src_payload~1_combout ),
	.src_payload2(\cmd_mux_014|src_payload~2_combout ),
	.src_payload3(\cmd_mux_014|src_payload~3_combout ),
	.src_payload4(\cmd_mux_014|src_payload~4_combout ),
	.src_payload5(\cmd_mux_014|src_payload~5_combout ),
	.src_payload6(\cmd_mux_014|src_payload~6_combout ),
	.src_payload7(\cmd_mux_014|src_payload~7_combout ),
	.src_data_105(\cmd_mux_014|src_data[105]~combout ),
	.src_data_106(\cmd_mux_014|src_data[106]~combout ),
	.src_data_107(\cmd_mux_014|src_data[107]~combout ),
	.src_data_108(\cmd_mux_014|src_data[108]~combout ),
	.src_data_109(\cmd_mux_014|src_data[109]~combout ),
	.src_data_110(\cmd_mux_014|src_data[110]~combout ),
	.src_data_111(\cmd_mux_014|src_data[111]~combout ),
	.src_data_112(\cmd_mux_014|src_data[112]~combout ),
	.src_data_113(\cmd_mux_014|src_data[113]~combout ),
	.src_data_114(\cmd_mux_014|src_data[114]~combout ),
	.src_data_115(\cmd_mux_014|src_data[115]~combout ),
	.src_data_116(\cmd_mux_014|src_data[116]~combout ),
	.src_data_86(\cmd_mux_014|src_data[86]~combout ),
	.Selector5(\hps_0_h2f_axi_master_agent|Selector5~1_combout ),
	.Selector12(\hps_0_h2f_axi_master_agent|Selector12~0_combout ),
	.out_data_1(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[1]~5_combout ),
	.src_data_80(\cmd_mux_014|src_data[80]~combout ),
	.out_data_0(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[0]~6_combout ),
	.Selector6(\hps_0_h2f_axi_master_agent|Selector6~0_combout ),
	.Selector13(\hps_0_h2f_axi_master_agent|Selector13~1_combout ),
	.src_data_79(\cmd_mux_014|src_data[79]~combout ),
	.clk_clk(clk_clk));

spw_babasu_altera_merlin_burst_adapter_10 tick_in_s1_burst_adapter(
	.h2f_ARADDR_0(h2f_ARADDR_0),
	.h2f_ARADDR_1(h2f_ARADDR_1),
	.h2f_ARADDR_2(h2f_ARADDR_2),
	.h2f_ARADDR_3(h2f_ARADDR_3),
	.h2f_ARLEN_0(h2f_ARLEN_0),
	.nxt_in_ready(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.in_ready_hold(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.stateST_COMP_TRANS(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.out_valid_reg(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.in_narrow_reg(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.in_byteen_reg_3(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ),
	.in_byteen_reg_2(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ),
	.in_byteen_reg_1(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ),
	.in_byteen_reg_0(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ),
	.in_data_reg_68(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ),
	.cp_ready(\tick_in_s1_agent|cp_ready~0_combout ),
	.stateST_UNCOMP_WR_SUBBURST(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.nxt_in_ready1(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.saved_grant_1(\cmd_mux_013|saved_grant[1]~q ),
	.Equal13(\router|Equal13~0_combout ),
	.saved_grant_0(\cmd_mux_013|saved_grant[0]~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.in_data_reg_0(in_data_reg_06),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_36),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_26),
	.Add2(\hps_0_h2f_axi_master_agent|Add2~0_combout ),
	.Add21(\hps_0_h2f_axi_master_agent|Add2~1_combout ),
	.Add22(\hps_0_h2f_axi_master_agent|Add2~2_combout ),
	.Add23(\hps_0_h2f_axi_master_agent|Add2~3_combout ),
	.Equal5(\router|Equal5~1_combout ),
	.write_cp_data_77(\hps_0_h2f_axi_master_agent|write_cp_data[77]~0_combout ),
	.write_cp_data_78(\hps_0_h2f_axi_master_agent|write_cp_data[78]~1_combout ),
	.write_cp_data_75(\hps_0_h2f_axi_master_agent|write_cp_data[75]~2_combout ),
	.write_cp_data_74(\hps_0_h2f_axi_master_agent|write_cp_data[74]~3_combout ),
	.write_cp_data_76(\hps_0_h2f_axi_master_agent|write_cp_data[76]~4_combout ),
	.WideNor0(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|WideNor0~0_combout ),
	.nxt_out_eop(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.src13_valid(\cmd_demux|src13_valid~1_combout ),
	.src_valid(\cmd_mux_013|src_valid~2_combout ),
	.cp_ready1(\tick_in_s1_agent|cp_ready~3_combout ),
	.in_data_reg_69(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.src_data_87(\cmd_mux_013|src_data[87]~combout ),
	.src_data_88(\cmd_mux_013|src_data[88]~combout ),
	.src_valid1(\cmd_mux_013|src_valid~3_combout ),
	.src_data_35(\cmd_mux_013|src_data[35]~combout ),
	.src_data_34(\cmd_mux_013|src_data[34]~combout ),
	.src_data_33(\cmd_mux_013|src_data[33]~combout ),
	.src_data_32(\cmd_mux_013|src_data[32]~combout ),
	.out_byte_cnt_reg_2(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_5(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_4(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_3(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_6(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.src_payload_0(\cmd_mux_013|src_payload[0]~combout ),
	.in_data_reg_105(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ),
	.in_data_reg_106(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ),
	.in_data_reg_107(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ),
	.in_data_reg_108(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ),
	.in_data_reg_109(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ),
	.in_data_reg_110(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ),
	.in_data_reg_111(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ),
	.in_data_reg_112(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ),
	.in_data_reg_113(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ),
	.in_data_reg_114(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ),
	.in_data_reg_115(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ),
	.in_data_reg_116(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ),
	.Selector3(\hps_0_h2f_axi_master_agent|Selector3~0_combout ),
	.Selector10(\hps_0_h2f_axi_master_agent|Selector10~1_combout ),
	.base_address_3(\hps_0_h2f_axi_master_agent|align_address_to_size|base_address[3]~0_combout ),
	.Selector4(\hps_0_h2f_axi_master_agent|Selector4~1_combout ),
	.Selector11(\hps_0_h2f_axi_master_agent|Selector11~1_combout ),
	.base_address_2(\hps_0_h2f_axi_master_agent|align_address_to_size|base_address[2]~1_combout ),
	.src_payload(\cmd_mux_013|src_payload~0_combout ),
	.src_data_82(\cmd_mux_013|src_data[82]~combout ),
	.src_data_81(\cmd_mux_013|src_data[81]~combout ),
	.src_data_105(\cmd_mux_013|src_data[105]~combout ),
	.src_data_106(\cmd_mux_013|src_data[106]~combout ),
	.src_data_107(\cmd_mux_013|src_data[107]~combout ),
	.src_data_108(\cmd_mux_013|src_data[108]~combout ),
	.src_data_109(\cmd_mux_013|src_data[109]~combout ),
	.src_data_110(\cmd_mux_013|src_data[110]~combout ),
	.src_data_111(\cmd_mux_013|src_data[111]~combout ),
	.src_data_112(\cmd_mux_013|src_data[112]~combout ),
	.src_data_113(\cmd_mux_013|src_data[113]~combout ),
	.src_data_114(\cmd_mux_013|src_data[114]~combout ),
	.src_data_115(\cmd_mux_013|src_data[115]~combout ),
	.src_data_116(\cmd_mux_013|src_data[116]~combout ),
	.src_data_86(\cmd_mux_013|src_data[86]~combout ),
	.Selector5(\hps_0_h2f_axi_master_agent|Selector5~1_combout ),
	.Selector12(\hps_0_h2f_axi_master_agent|Selector12~0_combout ),
	.out_data_1(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[1]~5_combout ),
	.src_data_80(\cmd_mux_013|src_data[80]~combout ),
	.out_data_0(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[0]~6_combout ),
	.Selector6(\hps_0_h2f_axi_master_agent|Selector6~0_combout ),
	.Selector13(\hps_0_h2f_axi_master_agent|Selector13~1_combout ),
	.src_data_79(\cmd_mux_013|src_data[79]~combout ),
	.clk_clk(clk_clk));

spw_babasu_altera_merlin_burst_adapter_1 currentstate_s1_burst_adapter(
	.h2f_ARADDR_0(h2f_ARADDR_0),
	.h2f_ARADDR_1(h2f_ARADDR_1),
	.h2f_ARADDR_2(h2f_ARADDR_2),
	.h2f_ARADDR_3(h2f_ARADDR_3),
	.h2f_ARBURST_0(h2f_ARBURST_0),
	.h2f_ARBURST_1(h2f_ARBURST_1),
	.h2f_ARID_0(h2f_ARID_0),
	.h2f_ARID_1(h2f_ARID_1),
	.h2f_ARID_2(h2f_ARID_2),
	.h2f_ARID_3(h2f_ARID_3),
	.h2f_ARID_4(h2f_ARID_4),
	.h2f_ARID_5(h2f_ARID_5),
	.h2f_ARID_6(h2f_ARID_6),
	.h2f_ARID_7(h2f_ARID_7),
	.h2f_ARID_8(h2f_ARID_8),
	.h2f_ARID_9(h2f_ARID_9),
	.h2f_ARID_10(h2f_ARID_10),
	.h2f_ARID_11(h2f_ARID_11),
	.h2f_ARLEN_0(h2f_ARLEN_0),
	.Add5(\hps_0_h2f_axi_master_agent|Add5~1_sumout ),
	.Add51(\hps_0_h2f_axi_master_agent|Add5~5_sumout ),
	.in_ready_hold(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.saved_grant_1(\cmd_mux_003|saved_grant[1]~q ),
	.stateST_COMP_TRANS(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.mem_used_1(\currentstate_s1_agent_rsp_fifo|mem_used[1]~q ),
	.in_data_reg_69(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.in_narrow_reg(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.cp_ready(\currentstate_s1_agent|cp_ready~0_combout ),
	.cp_ready1(\currentstate_s1_agent|cp_ready~1_combout ),
	.nxt_out_eop(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.out_valid_reg(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.stateST_UNCOMP_WR_SUBBURST(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.nxt_in_ready(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.Decoder1(\hps_0_h2f_axi_master_agent|Decoder1~0_combout ),
	.Add2(\hps_0_h2f_axi_master_agent|Add2~0_combout ),
	.Add21(\hps_0_h2f_axi_master_agent|Add2~1_combout ),
	.Add22(\hps_0_h2f_axi_master_agent|Add2~2_combout ),
	.Add23(\hps_0_h2f_axi_master_agent|Add2~3_combout ),
	.nxt_in_ready1(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.src_valid(\cmd_mux_003|src_valid~0_combout ),
	.out_byte_cnt_reg_2(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.cp_ready2(\currentstate_s1_agent|cp_ready~2_combout ),
	.out_uncomp_byte_cnt_reg_3(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_4(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_5(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_6(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.in_data_reg_105(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ),
	.in_data_reg_106(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ),
	.in_data_reg_107(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ),
	.in_data_reg_108(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ),
	.in_data_reg_109(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ),
	.in_data_reg_110(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ),
	.in_data_reg_111(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ),
	.in_data_reg_112(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ),
	.in_data_reg_113(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ),
	.in_data_reg_114(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ),
	.in_data_reg_115(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ),
	.in_data_reg_116(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ),
	.Selector10(\hps_0_h2f_axi_master_agent|Selector10~0_combout ),
	.Selector101(\hps_0_h2f_axi_master_agent|Selector10~1_combout ),
	.Selector11(\hps_0_h2f_axi_master_agent|Selector11~1_combout ),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_310),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_210),
	.Selector12(\hps_0_h2f_axi_master_agent|Selector12~0_combout ),
	.src_payload(\cmd_mux_003|src_payload~0_combout ),
	.src_payload1(\cmd_mux_003|src_payload~1_combout ),
	.src_payload2(\cmd_mux_003|src_payload~2_combout ),
	.Selector13(\hps_0_h2f_axi_master_agent|Selector13~1_combout ),
	.nxt_out_burstwrap_1(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_burstwrap[1]~0_combout ),
	.nxt_addr_2(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_addr[2]~2_combout ),
	.clk_clk(clk_clk));

spw_babasu_altera_merlin_burst_adapter autostart_s1_burst_adapter(
	.h2f_ARADDR_0(h2f_ARADDR_0),
	.h2f_ARADDR_1(h2f_ARADDR_1),
	.h2f_ARADDR_2(h2f_ARADDR_2),
	.h2f_ARADDR_3(h2f_ARADDR_3),
	.h2f_ARLEN_0(h2f_ARLEN_0),
	.nxt_in_ready(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.in_ready_hold(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.stateST_COMP_TRANS(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.out_valid_reg(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.in_narrow_reg(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.in_byteen_reg_3(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ),
	.in_byteen_reg_2(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ),
	.in_byteen_reg_1(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ),
	.in_byteen_reg_0(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ),
	.in_data_reg_68(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ),
	.cp_ready(\autostart_s1_agent|cp_ready~0_combout ),
	.stateST_UNCOMP_WR_SUBBURST(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.nxt_in_ready1(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.saved_grant_1(\cmd_mux_002|saved_grant[1]~q ),
	.Equal16(\router|Equal16~0_combout ),
	.saved_grant_0(\cmd_mux_002|saved_grant[0]~q ),
	.in_data_reg_0(in_data_reg_0),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_3),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_2),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.Add2(\hps_0_h2f_axi_master_agent|Add2~0_combout ),
	.Add21(\hps_0_h2f_axi_master_agent|Add2~1_combout ),
	.Add22(\hps_0_h2f_axi_master_agent|Add2~2_combout ),
	.Add23(\hps_0_h2f_axi_master_agent|Add2~3_combout ),
	.write_cp_data_77(\hps_0_h2f_axi_master_agent|write_cp_data[77]~0_combout ),
	.write_cp_data_78(\hps_0_h2f_axi_master_agent|write_cp_data[78]~1_combout ),
	.write_cp_data_75(\hps_0_h2f_axi_master_agent|write_cp_data[75]~2_combout ),
	.write_cp_data_74(\hps_0_h2f_axi_master_agent|write_cp_data[74]~3_combout ),
	.write_cp_data_76(\hps_0_h2f_axi_master_agent|write_cp_data[76]~4_combout ),
	.WideNor0(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|WideNor0~0_combout ),
	.Equal14(\router|Equal14~1_combout ),
	.nxt_out_eop(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.src2_valid(\cmd_demux|src2_valid~1_combout ),
	.src_valid(\cmd_mux_002|src_valid~0_combout ),
	.cp_ready1(\autostart_s1_agent|cp_ready~3_combout ),
	.in_data_reg_69(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.src_data_87(\cmd_mux_002|src_data[87]~combout ),
	.src_data_88(\cmd_mux_002|src_data[88]~combout ),
	.src_valid1(\cmd_mux_002|src_valid~1_combout ),
	.src_data_35(\cmd_mux_002|src_data[35]~combout ),
	.src_data_34(\cmd_mux_002|src_data[34]~combout ),
	.src_data_33(\cmd_mux_002|src_data[33]~combout ),
	.src_data_32(\cmd_mux_002|src_data[32]~combout ),
	.out_byte_cnt_reg_2(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_5(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_4(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_3(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_6(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.src_payload_0(\cmd_mux_002|src_payload[0]~combout ),
	.in_data_reg_105(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ),
	.in_data_reg_106(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ),
	.in_data_reg_107(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ),
	.in_data_reg_108(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ),
	.in_data_reg_109(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ),
	.in_data_reg_110(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ),
	.in_data_reg_111(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ),
	.in_data_reg_112(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ),
	.in_data_reg_113(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ),
	.in_data_reg_114(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ),
	.in_data_reg_115(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ),
	.in_data_reg_116(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ),
	.src_payload(\cmd_mux_002|src_payload~0_combout ),
	.Selector3(\hps_0_h2f_axi_master_agent|Selector3~0_combout ),
	.Selector10(\hps_0_h2f_axi_master_agent|Selector10~1_combout ),
	.src_data_82(\cmd_mux_002|src_data[82]~combout ),
	.base_address_3(\hps_0_h2f_axi_master_agent|align_address_to_size|base_address[3]~0_combout ),
	.Selector4(\hps_0_h2f_axi_master_agent|Selector4~1_combout ),
	.Selector11(\hps_0_h2f_axi_master_agent|Selector11~1_combout ),
	.src_data_81(\cmd_mux_002|src_data[81]~combout ),
	.base_address_2(\hps_0_h2f_axi_master_agent|align_address_to_size|base_address[2]~1_combout ),
	.src_data_105(\cmd_mux_002|src_data[105]~combout ),
	.src_data_106(\cmd_mux_002|src_data[106]~combout ),
	.src_data_107(\cmd_mux_002|src_data[107]~combout ),
	.src_data_108(\cmd_mux_002|src_data[108]~combout ),
	.src_data_109(\cmd_mux_002|src_data[109]~combout ),
	.src_data_110(\cmd_mux_002|src_data[110]~combout ),
	.src_data_111(\cmd_mux_002|src_data[111]~combout ),
	.src_data_112(\cmd_mux_002|src_data[112]~combout ),
	.src_data_113(\cmd_mux_002|src_data[113]~combout ),
	.src_data_114(\cmd_mux_002|src_data[114]~combout ),
	.src_data_115(\cmd_mux_002|src_data[115]~combout ),
	.src_data_116(\cmd_mux_002|src_data[116]~combout ),
	.src_data_86(\cmd_mux_002|src_data[86]~combout ),
	.Selector5(\hps_0_h2f_axi_master_agent|Selector5~1_combout ),
	.Selector12(\hps_0_h2f_axi_master_agent|Selector12~0_combout ),
	.src_data_80(\cmd_mux_002|src_data[80]~combout ),
	.out_data_1(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[1]~5_combout ),
	.out_data_0(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[0]~6_combout ),
	.Selector6(\hps_0_h2f_axi_master_agent|Selector6~0_combout ),
	.Selector13(\hps_0_h2f_axi_master_agent|Selector13~1_combout ),
	.src_data_79(\cmd_mux_002|src_data[79]~combout ),
	.clk_clk(clk_clk));

spw_babasu_altera_merlin_burst_adapter_5 link_disable_s1_burst_adapter(
	.h2f_ARADDR_0(h2f_ARADDR_0),
	.h2f_ARADDR_1(h2f_ARADDR_1),
	.h2f_ARADDR_2(h2f_ARADDR_2),
	.h2f_ARADDR_3(h2f_ARADDR_3),
	.h2f_ARLEN_0(h2f_ARLEN_0),
	.nxt_in_ready(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.in_ready_hold(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.stateST_COMP_TRANS(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.out_valid_reg(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.in_narrow_reg(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.in_byteen_reg_3(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ),
	.in_byteen_reg_2(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ),
	.in_byteen_reg_1(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ),
	.in_byteen_reg_0(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ),
	.in_data_reg_68(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ),
	.cp_ready(\link_disable_s1_agent|cp_ready~0_combout ),
	.stateST_UNCOMP_WR_SUBBURST(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.nxt_in_ready1(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.saved_grant_1(\cmd_mux_001|saved_grant[1]~q ),
	.Equal16(\router|Equal16~0_combout ),
	.saved_grant_0(\cmd_mux_001|saved_grant[0]~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.in_data_reg_0(in_data_reg_02),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_32),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_22),
	.Add2(\hps_0_h2f_axi_master_agent|Add2~0_combout ),
	.Add21(\hps_0_h2f_axi_master_agent|Add2~1_combout ),
	.Add22(\hps_0_h2f_axi_master_agent|Add2~2_combout ),
	.Add23(\hps_0_h2f_axi_master_agent|Add2~3_combout ),
	.nxt_out_eop(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.Equal5(\router|Equal5~1_combout ),
	.src1_valid(\cmd_demux|src1_valid~1_combout ),
	.src_valid(\cmd_mux_001|src_valid~0_combout ),
	.cp_ready1(\link_disable_s1_agent|cp_ready~3_combout ),
	.in_data_reg_69(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.src_data_87(\cmd_mux_001|src_data[87]~combout ),
	.src_data_88(\cmd_mux_001|src_data[88]~combout ),
	.src_valid1(\cmd_mux_001|src_valid~1_combout ),
	.src_data_35(\cmd_mux_001|src_data[35]~combout ),
	.src_data_34(\cmd_mux_001|src_data[34]~combout ),
	.src_data_33(\cmd_mux_001|src_data[33]~combout ),
	.src_data_32(\cmd_mux_001|src_data[32]~combout ),
	.out_byte_cnt_reg_2(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_3(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_4(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_5(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_6(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.src_payload_0(\cmd_mux_001|src_payload[0]~combout ),
	.write_cp_data_77(\hps_0_h2f_axi_master_agent|write_cp_data[77]~0_combout ),
	.write_cp_data_78(\hps_0_h2f_axi_master_agent|write_cp_data[78]~1_combout ),
	.write_cp_data_75(\hps_0_h2f_axi_master_agent|write_cp_data[75]~2_combout ),
	.write_cp_data_74(\hps_0_h2f_axi_master_agent|write_cp_data[74]~3_combout ),
	.write_cp_data_76(\hps_0_h2f_axi_master_agent|write_cp_data[76]~4_combout ),
	.WideNor0(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|WideNor0~0_combout ),
	.in_data_reg_105(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ),
	.in_data_reg_106(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ),
	.in_data_reg_107(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ),
	.in_data_reg_108(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ),
	.in_data_reg_109(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ),
	.in_data_reg_110(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ),
	.in_data_reg_111(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ),
	.in_data_reg_112(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ),
	.in_data_reg_113(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ),
	.in_data_reg_114(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ),
	.in_data_reg_115(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ),
	.in_data_reg_116(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ),
	.Selector3(\hps_0_h2f_axi_master_agent|Selector3~0_combout ),
	.Selector10(\hps_0_h2f_axi_master_agent|Selector10~1_combout ),
	.base_address_3(\hps_0_h2f_axi_master_agent|align_address_to_size|base_address[3]~0_combout ),
	.Selector4(\hps_0_h2f_axi_master_agent|Selector4~1_combout ),
	.Selector11(\hps_0_h2f_axi_master_agent|Selector11~1_combout ),
	.base_address_2(\hps_0_h2f_axi_master_agent|align_address_to_size|base_address[2]~1_combout ),
	.src_payload(\cmd_mux_001|src_payload~0_combout ),
	.src_data_82(\cmd_mux_001|src_data[82]~combout ),
	.src_data_81(\cmd_mux_001|src_data[81]~combout ),
	.src_data_105(\cmd_mux_001|src_data[105]~combout ),
	.src_data_106(\cmd_mux_001|src_data[106]~combout ),
	.src_data_107(\cmd_mux_001|src_data[107]~combout ),
	.src_data_108(\cmd_mux_001|src_data[108]~combout ),
	.src_data_109(\cmd_mux_001|src_data[109]~combout ),
	.src_data_110(\cmd_mux_001|src_data[110]~combout ),
	.src_data_111(\cmd_mux_001|src_data[111]~combout ),
	.src_data_112(\cmd_mux_001|src_data[112]~combout ),
	.src_data_113(\cmd_mux_001|src_data[113]~combout ),
	.src_data_114(\cmd_mux_001|src_data[114]~combout ),
	.src_data_115(\cmd_mux_001|src_data[115]~combout ),
	.src_data_116(\cmd_mux_001|src_data[116]~combout ),
	.src_data_86(\cmd_mux_001|src_data[86]~combout ),
	.Selector5(\hps_0_h2f_axi_master_agent|Selector5~1_combout ),
	.Selector12(\hps_0_h2f_axi_master_agent|Selector12~0_combout ),
	.out_data_1(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[1]~5_combout ),
	.src_data_80(\cmd_mux_001|src_data[80]~combout ),
	.out_data_0(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[0]~6_combout ),
	.Selector6(\hps_0_h2f_axi_master_agent|Selector6~0_combout ),
	.Selector13(\hps_0_h2f_axi_master_agent|Selector13~1_combout ),
	.src_data_79(\cmd_mux_001|src_data[79]~combout ),
	.clk_clk(clk_clk));

spw_babasu_altera_merlin_burst_adapter_6 link_start_s1_burst_adapter(
	.h2f_ARADDR_0(h2f_ARADDR_0),
	.h2f_ARADDR_1(h2f_ARADDR_1),
	.h2f_ARADDR_2(h2f_ARADDR_2),
	.h2f_ARADDR_3(h2f_ARADDR_3),
	.h2f_ARLEN_0(h2f_ARLEN_0),
	.nxt_in_ready(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~4_combout ),
	.in_ready_hold(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.saved_grant_1(\cmd_mux|saved_grant[1]~q ),
	.stateST_COMP_TRANS(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.out_valid_reg(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\link_start_s1_agent_rsp_fifo|mem_used[1]~q ),
	.in_narrow_reg(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.in_byteen_reg_3(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ),
	.in_byteen_reg_2(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ),
	.in_byteen_reg_1(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ),
	.in_byteen_reg_0(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ),
	.in_data_reg_68(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ),
	.cp_ready(\link_start_s1_agent|cp_ready~0_combout ),
	.stateST_UNCOMP_WR_SUBBURST(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.nxt_in_ready1(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.sop_enable(\hps_0_h2f_axi_master_agent|sop_enable~q ),
	.saved_grant_0(\cmd_mux|saved_grant[0]~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.in_data_reg_0(in_data_reg_03),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_33),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_23),
	.Add2(\hps_0_h2f_axi_master_agent|Add2~0_combout ),
	.Add21(\hps_0_h2f_axi_master_agent|Add2~1_combout ),
	.Add22(\hps_0_h2f_axi_master_agent|Add2~2_combout ),
	.Add23(\hps_0_h2f_axi_master_agent|Add2~3_combout ),
	.burst_bytecount_5(\hps_0_h2f_axi_master_agent|burst_bytecount[5]~q ),
	.write_cp_data_77(\hps_0_h2f_axi_master_agent|write_cp_data[77]~0_combout ),
	.burst_bytecount_6(\hps_0_h2f_axi_master_agent|burst_bytecount[6]~q ),
	.write_cp_data_78(\hps_0_h2f_axi_master_agent|write_cp_data[78]~1_combout ),
	.burst_bytecount_3(\hps_0_h2f_axi_master_agent|burst_bytecount[3]~q ),
	.write_cp_data_75(\hps_0_h2f_axi_master_agent|write_cp_data[75]~2_combout ),
	.burst_bytecount_2(\hps_0_h2f_axi_master_agent|burst_bytecount[2]~q ),
	.write_cp_data_74(\hps_0_h2f_axi_master_agent|write_cp_data[74]~3_combout ),
	.burst_bytecount_4(\hps_0_h2f_axi_master_agent|burst_bytecount[4]~q ),
	.write_cp_data_76(\hps_0_h2f_axi_master_agent|write_cp_data[76]~4_combout ),
	.WideNor0(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|WideNor0~0_combout ),
	.src0_valid(\cmd_demux|src0_valid~1_combout ),
	.src0_valid1(\cmd_demux_001|src0_valid~0_combout ),
	.nxt_in_ready2(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ),
	.src_valid(\cmd_mux|src_valid~0_combout ),
	.src_payload_0(\cmd_mux|src_payload[0]~combout ),
	.nxt_out_eop(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.cp_ready1(\link_start_s1_agent|cp_ready~2_combout ),
	.in_data_reg_69(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.src_data_87(\cmd_mux|src_data[87]~combout ),
	.src_data_88(\cmd_mux|src_data[88]~combout ),
	.src_data_35(\cmd_mux|src_data[35]~combout ),
	.src_data_34(\cmd_mux|src_data[34]~combout ),
	.src_data_33(\cmd_mux|src_data[33]~combout ),
	.src_data_32(\cmd_mux|src_data[32]~combout ),
	.out_byte_cnt_reg_2(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_3(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_4(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_5(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_6(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.in_data_reg_105(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ),
	.in_data_reg_106(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ),
	.in_data_reg_107(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ),
	.in_data_reg_108(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ),
	.in_data_reg_109(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ),
	.in_data_reg_110(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ),
	.in_data_reg_111(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ),
	.in_data_reg_112(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ),
	.in_data_reg_113(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ),
	.in_data_reg_114(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ),
	.in_data_reg_115(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ),
	.in_data_reg_116(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ),
	.Selector3(\hps_0_h2f_axi_master_agent|Selector3~0_combout ),
	.Selector10(\hps_0_h2f_axi_master_agent|Selector10~1_combout ),
	.base_address_3(\hps_0_h2f_axi_master_agent|align_address_to_size|base_address[3]~0_combout ),
	.Selector4(\hps_0_h2f_axi_master_agent|Selector4~1_combout ),
	.Selector11(\hps_0_h2f_axi_master_agent|Selector11~1_combout ),
	.base_address_2(\hps_0_h2f_axi_master_agent|align_address_to_size|base_address[2]~1_combout ),
	.src_payload(\cmd_mux|src_payload~0_combout ),
	.src_data_82(\cmd_mux|src_data[82]~combout ),
	.src_data_81(\cmd_mux|src_data[81]~combout ),
	.src_data_105(\cmd_mux|src_data[105]~combout ),
	.src_data_106(\cmd_mux|src_data[106]~combout ),
	.src_data_107(\cmd_mux|src_data[107]~combout ),
	.src_data_108(\cmd_mux|src_data[108]~combout ),
	.src_data_109(\cmd_mux|src_data[109]~combout ),
	.src_data_110(\cmd_mux|src_data[110]~combout ),
	.src_data_111(\cmd_mux|src_data[111]~combout ),
	.src_data_112(\cmd_mux|src_data[112]~combout ),
	.src_data_113(\cmd_mux|src_data[113]~combout ),
	.src_data_114(\cmd_mux|src_data[114]~combout ),
	.src_data_115(\cmd_mux|src_data[115]~combout ),
	.src_data_116(\cmd_mux|src_data[116]~combout ),
	.src_data_86(\cmd_mux|src_data[86]~combout ),
	.Selector5(\hps_0_h2f_axi_master_agent|Selector5~1_combout ),
	.Selector12(\hps_0_h2f_axi_master_agent|Selector12~0_combout ),
	.out_data_1(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[1]~5_combout ),
	.src_data_80(\cmd_mux|src_data[80]~combout ),
	.out_data_0(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[0]~6_combout ),
	.Selector6(\hps_0_h2f_axi_master_agent|Selector6~0_combout ),
	.Selector13(\hps_0_h2f_axi_master_agent|Selector13~1_combout ),
	.src_data_79(\cmd_mux|src_data[79]~combout ),
	.clk_clk(clk_clk));

spw_babasu_altera_merlin_traffic_limiter hps_0_h2f_axi_master_rd_limiter(
	.h2f_ARVALID_0(h2f_ARVALID_0),
	.h2f_RREADY_0(h2f_RREADY_0),
	.has_pending_responses1(\hps_0_h2f_axi_master_rd_limiter|has_pending_responses~q ),
	.cmd_sink_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\router_001|src_data[103]~3_combout ,\router_001|src_data[102]~0_combout ,\router_001|src_data[101]~2_combout ,\router_001|src_data[100]~1_combout ,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd}),
	.last_channel_6(\hps_0_h2f_axi_master_rd_limiter|last_channel[6]~q ),
	.cmd_sink_channel({\router_001|Equal16~0_combout ,\router_001|Equal15~0_combout ,\router_001|Equal14~0_combout ,\router_001|src_channel[13]~2_combout ,\cmd_mux_012|last_cycle~0_combout ,\cmd_mux_011|last_cycle~0_combout ,\router_001|Equal10~0_combout ,\router_001|Equal9~0_combout ,
\router_001|src_channel~0_combout ,\router_001|Equal7~0_combout ,\router_001|Equal6~0_combout ,\router_001|src_channel~5_combout ,\router_001|Equal4~0_combout ,\router_001|Equal3~0_combout ,\router_001|src_channel[2]~4_combout ,
\router_001|src_channel[1]~1_combout ,\router_001|src_channel[0]~3_combout }),
	.WideOr0(\cmd_demux_001|WideOr0~0_combout ),
	.WideOr01(\cmd_demux_001|WideOr0~1_combout ),
	.WideOr02(\cmd_demux_001|WideOr0~2_combout ),
	.WideOr03(\cmd_demux_001|WideOr0~6_combout ),
	.cmd_sink_ready(cmd_sink_ready),
	.src_payload(\rsp_mux_001|src_payload~0_combout ),
	.src_payload_0(\rsp_mux_001|src_payload[0]~6_combout ),
	.src_payload_01(\rsp_mux_001|src_payload[0]~13_combout ),
	.src_payload_02(\rsp_mux_001|src_payload[0]~19_combout ),
	.WideOr1(WideOr11),
	.reset(altera_reset_synchronizer_int_chain_out1),
	.last_channel_8(\hps_0_h2f_axi_master_rd_limiter|last_channel[8]~q ),
	.last_channel_11(\hps_0_h2f_axi_master_rd_limiter|last_channel[11]~q ),
	.last_channel_12(\hps_0_h2f_axi_master_rd_limiter|last_channel[12]~q ),
	.last_channel_1(\hps_0_h2f_axi_master_rd_limiter|last_channel[1]~q ),
	.last_channel_15(\hps_0_h2f_axi_master_rd_limiter|last_channel[15]~q ),
	.last_channel_16(\hps_0_h2f_axi_master_rd_limiter|last_channel[16]~q ),
	.last_channel_13(\hps_0_h2f_axi_master_rd_limiter|last_channel[13]~q ),
	.last_channel_14(\hps_0_h2f_axi_master_rd_limiter|last_channel[14]~q ),
	.last_channel_3(\hps_0_h2f_axi_master_rd_limiter|last_channel[3]~q ),
	.cmd_src_valid_5(\hps_0_h2f_axi_master_rd_limiter|cmd_src_valid[5]~0_combout ),
	.last_channel_9(\hps_0_h2f_axi_master_rd_limiter|last_channel[9]~q ),
	.last_channel_10(\hps_0_h2f_axi_master_rd_limiter|last_channel[10]~q ),
	.last_channel_0(\hps_0_h2f_axi_master_rd_limiter|last_channel[0]~q ),
	.last_channel_4(\hps_0_h2f_axi_master_rd_limiter|last_channel[4]~q ),
	.last_channel_7(\hps_0_h2f_axi_master_rd_limiter|last_channel[7]~q ),
	.last_channel_2(\hps_0_h2f_axi_master_rd_limiter|last_channel[2]~q ),
	.clk(clk_clk));

spw_babasu_altera_merlin_traffic_limiter_1 hps_0_h2f_axi_master_wr_limiter(
	.h2f_BREADY_0(h2f_BREADY_0),
	.h2f_WLAST_0(h2f_WLAST_0),
	.write_addr_data_both_valid(\hps_0_h2f_axi_master_agent|write_addr_data_both_valid~combout ),
	.has_pending_responses1(\hps_0_h2f_axi_master_wr_limiter|has_pending_responses~q ),
	.out_data_4(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[4]~2_combout ),
	.cmd_sink_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\router|src_data[103]~3_combout ,\router|src_data[102]~0_combout ,\router|src_data[101]~2_combout ,\router|src_data[100]~1_combout ,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.Equal5(\router|Equal5~0_combout ),
	.Equal14(\router|Equal14~0_combout ),
	.last_channel_6(\hps_0_h2f_axi_master_wr_limiter|last_channel[6]~q ),
	.WideOr0(\cmd_demux|WideOr0~0_combout ),
	.WideOr01(\cmd_demux|WideOr0~1_combout ),
	.WideOr02(\cmd_demux|WideOr0~2_combout ),
	.WideOr03(\cmd_demux|WideOr0~3_combout ),
	.WideOr04(\cmd_demux|WideOr0~4_combout ),
	.WideOr05(\cmd_demux|WideOr0~5_combout ),
	.nonposted_cmd_accepted(nonposted_cmd_accepted),
	.WideOr1(WideOr1),
	.nonposted_cmd_accepted1(nonposted_cmd_accepted1),
	.reset(altera_reset_synchronizer_int_chain_out1),
	.last_channel_1(\hps_0_h2f_axi_master_wr_limiter|last_channel[1]~q ),
	.last_channel_15(\hps_0_h2f_axi_master_wr_limiter|last_channel[15]~q ),
	.last_channel_16(\hps_0_h2f_axi_master_wr_limiter|last_channel[16]~q ),
	.last_channel_13(\hps_0_h2f_axi_master_wr_limiter|last_channel[13]~q ),
	.last_channel_14(\hps_0_h2f_axi_master_wr_limiter|last_channel[14]~q ),
	.last_channel_5(\hps_0_h2f_axi_master_wr_limiter|last_channel[5]~q ),
	.last_channel_9(\hps_0_h2f_axi_master_wr_limiter|last_channel[9]~q ),
	.last_channel_0(\hps_0_h2f_axi_master_wr_limiter|last_channel[0]~q ),
	.last_channel_2(\hps_0_h2f_axi_master_wr_limiter|last_channel[2]~q ),
	.src_payload(\rsp_mux|src_payload~0_combout ),
	.src_payload1(\rsp_mux|src_payload~1_combout ),
	.src_payload_0(\rsp_mux|src_payload[0]~8_combout ),
	.src_payload_01(\rsp_mux|src_payload[0]~9_combout ),
	.cmd_sink_channel({\router|Equal16~2_combout ,\router|Equal15~2_combout ,\router|Equal14~2_combout ,\router|Equal13~1_combout ,gnd,gnd,gnd,\router|Equal9~1_combout ,gnd,gnd,\router|Equal6~0_combout ,\router|Equal5~2_combout ,gnd,gnd,\router|Equal2~0_combout ,\router|src_channel~0_combout ,
\router|src_channel[0]~1_combout }),
	.clk(clk_clk));

spw_babasu_altera_merlin_slave_agent_9 spill_enable_s1_agent(
	.waitrequest_reset_override(\autostart_s1_translator|waitrequest_reset_override~q ),
	.stateST_COMP_TRANS(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.out_valid_reg(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\spill_enable_s1_agent_rsp_fifo|mem_used[1]~q ),
	.in_narrow_reg(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.in_byteen_reg_3(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ),
	.in_byteen_reg_2(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ),
	.in_byteen_reg_1(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ),
	.in_byteen_reg_0(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ),
	.WideOr0(\spill_enable_s1_agent|WideOr0~0_combout ),
	.wait_latency_counter_1(wait_latency_counter_12),
	.wait_latency_counter_0(wait_latency_counter_02),
	.in_data_reg_68(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ),
	.cp_ready(\spill_enable_s1_agent|cp_ready~0_combout ),
	.read_latency_shift_reg_0(\spill_enable_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\spill_enable_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_129_0(\spill_enable_s1_agent_rsp_fifo|mem[0][129]~q ),
	.mem_used_01(\spill_enable_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_66_0(\spill_enable_s1_agent_rsp_fifo|mem[0][66]~q ),
	.comb(\spill_enable_s1_agent|comb~0_combout ),
	.last_packet_beat(\spill_enable_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.mem_78_0(\spill_enable_s1_agent_rsp_fifo|mem[0][78]~q ),
	.mem_77_0(\spill_enable_s1_agent_rsp_fifo|mem[0][77]~q ),
	.mem_76_0(\spill_enable_s1_agent_rsp_fifo|mem[0][76]~q ),
	.mem_75_0(\spill_enable_s1_agent_rsp_fifo|mem[0][75]~q ),
	.mem_74_0(\spill_enable_s1_agent_rsp_fifo|mem[0][74]~q ),
	.last_packet_beat1(\spill_enable_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.m0_write1(m0_write5),
	.nxt_out_eop(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.cp_ready1(\spill_enable_s1_agent|cp_ready~1_combout ),
	.cp_ready2(\spill_enable_s1_agent|cp_ready~2_combout ),
	.last_packet_beat2(\spill_enable_s1_agent|uncompressor|last_packet_beat~2_combout ),
	.WideOr01(\rsp_demux_016|WideOr0~0_combout ),
	.read(\spill_enable_s1_agent_rsp_fifo|read~0_combout ),
	.cp_ready3(\spill_enable_s1_agent|cp_ready~3_combout ),
	.in_data_reg_69(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.rf_source_valid(\spill_enable_s1_agent|rf_source_valid~0_combout ),
	.rf_sink_ready(\spill_enable_s1_agent|uncompressor|sink_ready~0_combout ),
	.clk_clk(clk_clk));

spw_babasu_altera_avalon_sc_fifo_28 tx_clk_div_s1_agent_rdata_fifo(
	.read_latency_shift_reg_0(\tx_clk_div_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\tx_clk_div_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_129_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][129]~q ),
	.mem_used_01(\tx_clk_div_s1_agent_rsp_fifo|mem_used[0]~q ),
	.av_readdata_pre_0(\tx_clk_div_s1_translator|av_readdata_pre[0]~q ),
	.always4(\tx_clk_div_s1_agent_rdata_fifo|always4~0_combout ),
	.mem_0_0(\tx_clk_div_s1_agent_rdata_fifo|mem[0][0]~q ),
	.av_readdata_pre_1(\tx_clk_div_s1_translator|av_readdata_pre[1]~q ),
	.mem_1_0(\tx_clk_div_s1_agent_rdata_fifo|mem[0][1]~q ),
	.av_readdata_pre_2(\tx_clk_div_s1_translator|av_readdata_pre[2]~q ),
	.mem_2_0(\tx_clk_div_s1_agent_rdata_fifo|mem[0][2]~q ),
	.av_readdata_pre_3(\tx_clk_div_s1_translator|av_readdata_pre[3]~q ),
	.mem_3_0(\tx_clk_div_s1_agent_rdata_fifo|mem[0][3]~q ),
	.av_readdata_pre_4(\tx_clk_div_s1_translator|av_readdata_pre[4]~q ),
	.mem_4_0(\tx_clk_div_s1_agent_rdata_fifo|mem[0][4]~q ),
	.av_readdata_pre_5(\tx_clk_div_s1_translator|av_readdata_pre[5]~q ),
	.mem_5_0(\tx_clk_div_s1_agent_rdata_fifo|mem[0][5]~q ),
	.av_readdata_pre_6(\tx_clk_div_s1_translator|av_readdata_pre[6]~q ),
	.mem_6_0(\tx_clk_div_s1_agent_rdata_fifo|mem[0][6]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.WideOr0(\rsp_demux_015|WideOr0~0_combout ),
	.clk(clk_clk));

spw_babasu_altera_avalon_sc_fifo_29 tx_clk_div_s1_agent_rsp_fifo(
	.out_valid_reg(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\tx_clk_div_s1_agent_rsp_fifo|mem_used[1]~q ),
	.WideOr0(\tx_clk_div_s1_agent|WideOr0~0_combout ),
	.in_data_reg_68(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ),
	.stateST_UNCOMP_WR_SUBBURST(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.mem_129_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][129]~q ),
	.mem_used_0(\tx_clk_div_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_68_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][68]~q ),
	.mem_66_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][66]~q ),
	.comb(\tx_clk_div_s1_agent|comb~0_combout ),
	.mem_130_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][130]~q ),
	.mem_78_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][78]~q ),
	.mem_77_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][77]~q ),
	.mem_76_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][76]~q ),
	.mem_75_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][75]~q ),
	.mem_74_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][74]~q ),
	.mem_105_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][105]~q ),
	.mem_106_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][106]~q ),
	.mem_107_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][107]~q ),
	.mem_108_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][108]~q ),
	.mem_109_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][109]~q ),
	.mem_110_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][110]~q ),
	.mem_111_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][111]~q ),
	.mem_112_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_113_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][113]~q ),
	.mem_114_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][114]~q ),
	.mem_115_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][115]~q ),
	.mem_116_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][116]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.nxt_out_eop(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.last_packet_beat(\tx_clk_div_s1_agent|uncompressor|last_packet_beat~2_combout ),
	.WideOr01(\rsp_demux_015|WideOr0~0_combout ),
	.read(\tx_clk_div_s1_agent_rsp_fifo|read~0_combout ),
	.cp_ready(\tx_clk_div_s1_agent|cp_ready~4_combout ),
	.in_data_reg_69(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.rf_source_valid(\tx_clk_div_s1_agent|rf_source_valid~0_combout ),
	.out_byte_cnt_reg_2(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_4(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_3(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_5(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_6(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.sink_ready(\tx_clk_div_s1_agent|uncompressor|sink_ready~0_combout ),
	.in_data_reg_105(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ),
	.in_data_reg_106(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ),
	.in_data_reg_107(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ),
	.in_data_reg_108(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ),
	.in_data_reg_109(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ),
	.in_data_reg_110(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ),
	.in_data_reg_111(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ),
	.in_data_reg_112(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ),
	.in_data_reg_113(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ),
	.in_data_reg_114(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ),
	.in_data_reg_115(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ),
	.in_data_reg_116(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ),
	.clk(clk_clk));

spw_babasu_altera_merlin_slave_agent_14 tx_clk_div_s1_agent(
	.waitrequest_reset_override(\autostart_s1_translator|waitrequest_reset_override~q ),
	.stateST_COMP_TRANS(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.out_valid_reg(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\tx_clk_div_s1_agent_rsp_fifo|mem_used[1]~q ),
	.in_narrow_reg(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.in_byteen_reg_3(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ),
	.in_byteen_reg_2(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ),
	.in_byteen_reg_1(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ),
	.in_byteen_reg_0(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ),
	.WideOr0(\tx_clk_div_s1_agent|WideOr0~0_combout ),
	.wait_latency_counter_1(wait_latency_counter_11),
	.wait_latency_counter_0(wait_latency_counter_01),
	.in_data_reg_68(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ),
	.cp_ready(\tx_clk_div_s1_agent|cp_ready~0_combout ),
	.read_latency_shift_reg_0(\tx_clk_div_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\tx_clk_div_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_129_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][129]~q ),
	.mem_used_01(\tx_clk_div_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_66_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][66]~q ),
	.comb(\tx_clk_div_s1_agent|comb~0_combout ),
	.last_packet_beat(\tx_clk_div_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.mem_78_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][78]~q ),
	.mem_77_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][77]~q ),
	.mem_76_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][76]~q ),
	.mem_75_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][75]~q ),
	.mem_74_0(\tx_clk_div_s1_agent_rsp_fifo|mem[0][74]~q ),
	.last_packet_beat1(\tx_clk_div_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.m0_write1(m0_write8),
	.nxt_out_eop(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.cp_ready1(\tx_clk_div_s1_agent|cp_ready~3_combout ),
	.last_packet_beat2(\tx_clk_div_s1_agent|uncompressor|last_packet_beat~2_combout ),
	.WideOr01(\rsp_demux_015|WideOr0~0_combout ),
	.read(\tx_clk_div_s1_agent_rsp_fifo|read~0_combout ),
	.cp_ready2(\tx_clk_div_s1_agent|cp_ready~4_combout ),
	.in_data_reg_69(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.rf_source_valid(\tx_clk_div_s1_agent|rf_source_valid~0_combout ),
	.rf_sink_ready(\tx_clk_div_s1_agent|uncompressor|sink_ready~0_combout ),
	.clk_clk(clk_clk));

spw_babasu_altera_avalon_sc_fifo_24 time_in_s1_agent_rdata_fifo(
	.read_latency_shift_reg_0(\time_in_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\time_in_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_129_0(\time_in_s1_agent_rsp_fifo|mem[0][129]~q ),
	.mem_used_01(\time_in_s1_agent_rsp_fifo|mem_used[0]~q ),
	.av_readdata_pre_0(\time_in_s1_translator|av_readdata_pre[0]~q ),
	.always4(\time_in_s1_agent_rdata_fifo|always4~0_combout ),
	.mem_0_0(\time_in_s1_agent_rdata_fifo|mem[0][0]~q ),
	.av_readdata_pre_1(\time_in_s1_translator|av_readdata_pre[1]~q ),
	.mem_1_0(\time_in_s1_agent_rdata_fifo|mem[0][1]~q ),
	.av_readdata_pre_2(\time_in_s1_translator|av_readdata_pre[2]~q ),
	.mem_2_0(\time_in_s1_agent_rdata_fifo|mem[0][2]~q ),
	.av_readdata_pre_3(\time_in_s1_translator|av_readdata_pre[3]~q ),
	.mem_3_0(\time_in_s1_agent_rdata_fifo|mem[0][3]~q ),
	.av_readdata_pre_4(\time_in_s1_translator|av_readdata_pre[4]~q ),
	.mem_4_0(\time_in_s1_agent_rdata_fifo|mem[0][4]~q ),
	.av_readdata_pre_5(\time_in_s1_translator|av_readdata_pre[5]~q ),
	.mem_5_0(\time_in_s1_agent_rdata_fifo|mem[0][5]~q ),
	.av_readdata_pre_6(\time_in_s1_translator|av_readdata_pre[6]~q ),
	.mem_6_0(\time_in_s1_agent_rdata_fifo|mem[0][6]~q ),
	.av_readdata_pre_7(\time_in_s1_translator|av_readdata_pre[7]~q ),
	.mem_7_0(\time_in_s1_agent_rdata_fifo|mem[0][7]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.WideOr0(\rsp_demux_014|WideOr0~0_combout ),
	.clk(clk_clk));

spw_babasu_altera_avalon_sc_fifo_25 time_in_s1_agent_rsp_fifo(
	.out_valid_reg(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\time_in_s1_agent_rsp_fifo|mem_used[1]~q ),
	.WideOr0(\time_in_s1_agent|WideOr0~0_combout ),
	.in_data_reg_68(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ),
	.stateST_UNCOMP_WR_SUBBURST(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.mem_129_0(\time_in_s1_agent_rsp_fifo|mem[0][129]~q ),
	.mem_used_0(\time_in_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_68_0(\time_in_s1_agent_rsp_fifo|mem[0][68]~q ),
	.mem_66_0(\time_in_s1_agent_rsp_fifo|mem[0][66]~q ),
	.comb(\time_in_s1_agent|comb~0_combout ),
	.mem_130_0(\time_in_s1_agent_rsp_fifo|mem[0][130]~q ),
	.mem_78_0(\time_in_s1_agent_rsp_fifo|mem[0][78]~q ),
	.mem_77_0(\time_in_s1_agent_rsp_fifo|mem[0][77]~q ),
	.mem_76_0(\time_in_s1_agent_rsp_fifo|mem[0][76]~q ),
	.mem_75_0(\time_in_s1_agent_rsp_fifo|mem[0][75]~q ),
	.mem_74_0(\time_in_s1_agent_rsp_fifo|mem[0][74]~q ),
	.mem_105_0(\time_in_s1_agent_rsp_fifo|mem[0][105]~q ),
	.mem_106_0(\time_in_s1_agent_rsp_fifo|mem[0][106]~q ),
	.mem_107_0(\time_in_s1_agent_rsp_fifo|mem[0][107]~q ),
	.mem_108_0(\time_in_s1_agent_rsp_fifo|mem[0][108]~q ),
	.mem_109_0(\time_in_s1_agent_rsp_fifo|mem[0][109]~q ),
	.mem_110_0(\time_in_s1_agent_rsp_fifo|mem[0][110]~q ),
	.mem_111_0(\time_in_s1_agent_rsp_fifo|mem[0][111]~q ),
	.mem_112_0(\time_in_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_113_0(\time_in_s1_agent_rsp_fifo|mem[0][113]~q ),
	.mem_114_0(\time_in_s1_agent_rsp_fifo|mem[0][114]~q ),
	.mem_115_0(\time_in_s1_agent_rsp_fifo|mem[0][115]~q ),
	.mem_116_0(\time_in_s1_agent_rsp_fifo|mem[0][116]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.nxt_out_eop(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.last_packet_beat(\time_in_s1_agent|uncompressor|last_packet_beat~2_combout ),
	.WideOr01(\rsp_demux_014|WideOr0~0_combout ),
	.read(\time_in_s1_agent_rsp_fifo|read~0_combout ),
	.cp_ready(\time_in_s1_agent|cp_ready~4_combout ),
	.in_data_reg_69(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.rf_source_valid(\time_in_s1_agent|rf_source_valid~0_combout ),
	.out_byte_cnt_reg_2(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_5(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_4(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_3(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_6(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.rp_valid(\time_in_s1_agent|rp_valid~combout ),
	.in_data_reg_105(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ),
	.in_data_reg_106(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ),
	.in_data_reg_107(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ),
	.in_data_reg_108(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ),
	.in_data_reg_109(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ),
	.in_data_reg_110(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ),
	.in_data_reg_111(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ),
	.in_data_reg_112(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ),
	.in_data_reg_113(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ),
	.in_data_reg_114(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ),
	.in_data_reg_115(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ),
	.in_data_reg_116(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ),
	.clk(clk_clk));

spw_babasu_altera_merlin_slave_agent_12 time_in_s1_agent(
	.waitrequest_reset_override(\autostart_s1_translator|waitrequest_reset_override~q ),
	.stateST_COMP_TRANS(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.out_valid_reg(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\time_in_s1_agent_rsp_fifo|mem_used[1]~q ),
	.in_narrow_reg(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.in_byteen_reg_3(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ),
	.in_byteen_reg_2(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ),
	.in_byteen_reg_1(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ),
	.in_byteen_reg_0(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ),
	.WideOr0(\time_in_s1_agent|WideOr0~0_combout ),
	.wait_latency_counter_1(wait_latency_counter_14),
	.wait_latency_counter_0(wait_latency_counter_04),
	.in_data_reg_68(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ),
	.cp_ready(\time_in_s1_agent|cp_ready~0_combout ),
	.read_latency_shift_reg_0(\time_in_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\time_in_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_129_0(\time_in_s1_agent_rsp_fifo|mem[0][129]~q ),
	.mem_used_01(\time_in_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_66_0(\time_in_s1_agent_rsp_fifo|mem[0][66]~q ),
	.comb(\time_in_s1_agent|comb~0_combout ),
	.last_packet_beat(\time_in_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.mem_78_0(\time_in_s1_agent_rsp_fifo|mem[0][78]~q ),
	.mem_77_0(\time_in_s1_agent_rsp_fifo|mem[0][77]~q ),
	.mem_76_0(\time_in_s1_agent_rsp_fifo|mem[0][76]~q ),
	.mem_75_0(\time_in_s1_agent_rsp_fifo|mem[0][75]~q ),
	.mem_74_0(\time_in_s1_agent_rsp_fifo|mem[0][74]~q ),
	.last_packet_beat1(\time_in_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.m0_write1(m0_write7),
	.nxt_out_eop(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.cp_ready1(\time_in_s1_agent|cp_ready~3_combout ),
	.last_packet_beat2(\time_in_s1_agent|uncompressor|last_packet_beat~2_combout ),
	.read(\time_in_s1_agent_rsp_fifo|read~0_combout ),
	.cp_ready2(\time_in_s1_agent|cp_ready~4_combout ),
	.in_data_reg_69(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.rf_source_valid(\time_in_s1_agent|rf_source_valid~0_combout ),
	.rp_valid1(\time_in_s1_agent|rp_valid~combout ),
	.clk_clk(clk_clk));

spw_babasu_altera_avalon_sc_fifo_20 tick_in_s1_agent_rdata_fifo(
	.read_latency_shift_reg_0(\tick_in_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\tick_in_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_129_0(\tick_in_s1_agent_rsp_fifo|mem[0][129]~q ),
	.mem_used_01(\tick_in_s1_agent_rsp_fifo|mem_used[0]~q ),
	.av_readdata_pre_0(\tick_in_s1_translator|av_readdata_pre[0]~q ),
	.mem_0_0(\tick_in_s1_agent_rdata_fifo|mem[0][0]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.WideOr0(\rsp_demux_013|WideOr0~0_combout ),
	.clk(clk_clk));

spw_babasu_altera_avalon_sc_fifo_21 tick_in_s1_agent_rsp_fifo(
	.out_valid_reg(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\tick_in_s1_agent_rsp_fifo|mem_used[1]~q ),
	.WideOr0(\tick_in_s1_agent|WideOr0~0_combout ),
	.in_data_reg_68(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ),
	.stateST_UNCOMP_WR_SUBBURST(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.mem_129_0(\tick_in_s1_agent_rsp_fifo|mem[0][129]~q ),
	.mem_used_0(\tick_in_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_68_0(\tick_in_s1_agent_rsp_fifo|mem[0][68]~q ),
	.mem_66_0(\tick_in_s1_agent_rsp_fifo|mem[0][66]~q ),
	.comb(\tick_in_s1_agent|comb~0_combout ),
	.mem_130_0(\tick_in_s1_agent_rsp_fifo|mem[0][130]~q ),
	.mem_78_0(\tick_in_s1_agent_rsp_fifo|mem[0][78]~q ),
	.mem_77_0(\tick_in_s1_agent_rsp_fifo|mem[0][77]~q ),
	.mem_76_0(\tick_in_s1_agent_rsp_fifo|mem[0][76]~q ),
	.mem_75_0(\tick_in_s1_agent_rsp_fifo|mem[0][75]~q ),
	.mem_74_0(\tick_in_s1_agent_rsp_fifo|mem[0][74]~q ),
	.mem_105_0(\tick_in_s1_agent_rsp_fifo|mem[0][105]~q ),
	.mem_106_0(\tick_in_s1_agent_rsp_fifo|mem[0][106]~q ),
	.mem_107_0(\tick_in_s1_agent_rsp_fifo|mem[0][107]~q ),
	.mem_108_0(\tick_in_s1_agent_rsp_fifo|mem[0][108]~q ),
	.mem_109_0(\tick_in_s1_agent_rsp_fifo|mem[0][109]~q ),
	.mem_110_0(\tick_in_s1_agent_rsp_fifo|mem[0][110]~q ),
	.mem_111_0(\tick_in_s1_agent_rsp_fifo|mem[0][111]~q ),
	.mem_112_0(\tick_in_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_113_0(\tick_in_s1_agent_rsp_fifo|mem[0][113]~q ),
	.mem_114_0(\tick_in_s1_agent_rsp_fifo|mem[0][114]~q ),
	.mem_115_0(\tick_in_s1_agent_rsp_fifo|mem[0][115]~q ),
	.mem_116_0(\tick_in_s1_agent_rsp_fifo|mem[0][116]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.nxt_out_eop(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.last_packet_beat(\tick_in_s1_agent|uncompressor|last_packet_beat~2_combout ),
	.WideOr01(\rsp_demux_013|WideOr0~0_combout ),
	.read(\tick_in_s1_agent_rsp_fifo|read~0_combout ),
	.cp_ready(\tick_in_s1_agent|cp_ready~4_combout ),
	.in_data_reg_69(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.rf_source_valid(\tick_in_s1_agent|rf_source_valid~0_combout ),
	.out_byte_cnt_reg_2(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_5(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_4(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_3(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_6(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.rp_valid(\tick_in_s1_agent|rp_valid~combout ),
	.in_data_reg_105(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ),
	.in_data_reg_106(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ),
	.in_data_reg_107(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ),
	.in_data_reg_108(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ),
	.in_data_reg_109(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ),
	.in_data_reg_110(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ),
	.in_data_reg_111(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ),
	.in_data_reg_112(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ),
	.in_data_reg_113(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ),
	.in_data_reg_114(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ),
	.in_data_reg_115(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ),
	.in_data_reg_116(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ),
	.clk(clk_clk));

spw_babasu_altera_merlin_slave_agent_10 tick_in_s1_agent(
	.waitrequest_reset_override(\autostart_s1_translator|waitrequest_reset_override~q ),
	.stateST_COMP_TRANS(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.out_valid_reg(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\tick_in_s1_agent_rsp_fifo|mem_used[1]~q ),
	.in_narrow_reg(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.in_byteen_reg_3(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ),
	.in_byteen_reg_2(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ),
	.in_byteen_reg_1(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ),
	.in_byteen_reg_0(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ),
	.WideOr0(\tick_in_s1_agent|WideOr0~0_combout ),
	.wait_latency_counter_1(wait_latency_counter_13),
	.wait_latency_counter_0(wait_latency_counter_03),
	.in_data_reg_68(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ),
	.cp_ready(\tick_in_s1_agent|cp_ready~0_combout ),
	.read_latency_shift_reg_0(\tick_in_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\tick_in_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_129_0(\tick_in_s1_agent_rsp_fifo|mem[0][129]~q ),
	.mem_used_01(\tick_in_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_66_0(\tick_in_s1_agent_rsp_fifo|mem[0][66]~q ),
	.comb(\tick_in_s1_agent|comb~0_combout ),
	.last_packet_beat(\tick_in_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.mem_78_0(\tick_in_s1_agent_rsp_fifo|mem[0][78]~q ),
	.mem_77_0(\tick_in_s1_agent_rsp_fifo|mem[0][77]~q ),
	.mem_76_0(\tick_in_s1_agent_rsp_fifo|mem[0][76]~q ),
	.mem_75_0(\tick_in_s1_agent_rsp_fifo|mem[0][75]~q ),
	.mem_74_0(\tick_in_s1_agent_rsp_fifo|mem[0][74]~q ),
	.last_packet_beat1(\tick_in_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.m0_write1(m0_write6),
	.nxt_out_eop(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.cp_ready1(\tick_in_s1_agent|cp_ready~3_combout ),
	.last_packet_beat2(\tick_in_s1_agent|uncompressor|last_packet_beat~2_combout ),
	.read(\tick_in_s1_agent_rsp_fifo|read~0_combout ),
	.cp_ready2(\tick_in_s1_agent|cp_ready~4_combout ),
	.in_data_reg_69(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.rf_source_valid(\tick_in_s1_agent|rf_source_valid~0_combout ),
	.rp_valid1(\tick_in_s1_agent|rp_valid~combout ),
	.clk_clk(clk_clk));

spw_babasu_altera_avalon_sc_fifo_26 time_out_s1_agent_rdata_fifo(
	.h2f_RREADY_0(h2f_RREADY_0),
	.read_latency_shift_reg_0(\time_out_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\time_out_s1_agent_rdata_fifo|mem_used[0]~q ),
	.empty1(\time_out_s1_agent_rdata_fifo|empty~combout ),
	.mem_0_0(\time_out_s1_agent_rdata_fifo|mem[0][0]~q ),
	.av_readdata_pre_0(\time_out_s1_translator|av_readdata_pre[0]~q ),
	.mem_1_0(\time_out_s1_agent_rdata_fifo|mem[0][1]~q ),
	.av_readdata_pre_1(\time_out_s1_translator|av_readdata_pre[1]~q ),
	.mem_2_0(\time_out_s1_agent_rdata_fifo|mem[0][2]~q ),
	.av_readdata_pre_2(\time_out_s1_translator|av_readdata_pre[2]~q ),
	.mem_3_0(\time_out_s1_agent_rdata_fifo|mem[0][3]~q ),
	.av_readdata_pre_3(\time_out_s1_translator|av_readdata_pre[3]~q ),
	.mem_4_0(\time_out_s1_agent_rdata_fifo|mem[0][4]~q ),
	.av_readdata_pre_4(\time_out_s1_translator|av_readdata_pre[4]~q ),
	.mem_5_0(\time_out_s1_agent_rdata_fifo|mem[0][5]~q ),
	.av_readdata_pre_5(\time_out_s1_translator|av_readdata_pre[5]~q ),
	.mem_6_0(\time_out_s1_agent_rdata_fifo|mem[0][6]~q ),
	.av_readdata_pre_6(\time_out_s1_translator|av_readdata_pre[6]~q ),
	.mem_7_0(\time_out_s1_agent_rdata_fifo|mem[0][7]~q ),
	.av_readdata_pre_7(\time_out_s1_translator|av_readdata_pre[7]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.clk(clk_clk));

spw_babasu_spw_babasu_mm_interconnect_0_router_1 router_001(
	.h2f_ARADDR_4(h2f_ARADDR_4),
	.h2f_ARADDR_5(h2f_ARADDR_5),
	.h2f_ARADDR_6(h2f_ARADDR_6),
	.h2f_ARADDR_7(h2f_ARADDR_7),
	.h2f_ARADDR_8(h2f_ARADDR_8),
	.src_data_102(\router_001|src_data[102]~0_combout ),
	.Equal6(\router_001|Equal6~0_combout ),
	.src_data_100(\router_001|src_data[100]~1_combout ),
	.src_data_101(\router_001|src_data[101]~2_combout ),
	.src_data_103(\router_001|src_data[103]~3_combout ),
	.src_channel(\router_001|src_channel~0_combout ),
	.src_channel_1(\router_001|src_channel[1]~1_combout ),
	.Equal15(\router_001|Equal15~0_combout ),
	.Equal16(\router_001|Equal16~0_combout ),
	.src_channel_13(\router_001|src_channel[13]~2_combout ),
	.Equal14(\router_001|Equal14~0_combout ),
	.Equal3(\router_001|Equal3~0_combout ),
	.Equal10(\router_001|Equal10~0_combout ),
	.src_channel_0(\router_001|src_channel[0]~3_combout ),
	.Equal9(\router_001|Equal9~0_combout ),
	.Equal4(\router_001|Equal4~0_combout ),
	.Equal7(\router_001|Equal7~0_combout ),
	.src_channel_2(\router_001|src_channel[2]~4_combout ),
	.src_channel1(\router_001|src_channel~5_combout ));

spw_babasu_spw_babasu_mm_interconnect_0_router router(
	.h2f_AWADDR_4(h2f_AWADDR_4),
	.h2f_AWADDR_5(h2f_AWADDR_5),
	.h2f_AWADDR_6(h2f_AWADDR_6),
	.h2f_AWADDR_7(h2f_AWADDR_7),
	.h2f_AWADDR_8(h2f_AWADDR_8),
	.address_burst_8(\hps_0_h2f_axi_master_agent|align_address_to_size|address_burst[8]~q ),
	.address_burst_7(\hps_0_h2f_axi_master_agent|align_address_to_size|address_burst[7]~q ),
	.address_burst_6(\hps_0_h2f_axi_master_agent|align_address_to_size|address_burst[6]~q ),
	.sop_enable(\hps_0_h2f_axi_master_agent|sop_enable~q ),
	.out_data_8(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[8]~0_combout ),
	.address_burst_5(\hps_0_h2f_axi_master_agent|align_address_to_size|address_burst[5]~q ),
	.out_data_5(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[5]~1_combout ),
	.address_burst_4(\hps_0_h2f_axi_master_agent|align_address_to_size|address_burst[4]~q ),
	.out_data_4(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[4]~2_combout ),
	.out_data_7(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[7]~3_combout ),
	.out_data_6(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[6]~4_combout ),
	.src_data_102(\router|src_data[102]~0_combout ),
	.Equal5(\router|Equal5~0_combout ),
	.Equal14(\router|Equal14~0_combout ),
	.src_data_100(\router|src_data[100]~1_combout ),
	.src_data_101(\router|src_data[101]~2_combout ),
	.Equal16(\router|Equal16~0_combout ),
	.Equal13(\router|Equal13~0_combout ),
	.src_data_103(\router|src_data[103]~3_combout ),
	.Equal15(\router|Equal15~0_combout ),
	.Equal161(\router|Equal16~1_combout ),
	.Equal9(\router|Equal9~0_combout ),
	.Equal51(\router|Equal5~1_combout ),
	.Equal151(\router|Equal15~1_combout ),
	.Equal141(\router|Equal14~1_combout ),
	.Equal6(\router|Equal6~0_combout ),
	.src_channel(\router|src_channel~0_combout ),
	.Equal152(\router|Equal15~2_combout ),
	.Equal162(\router|Equal16~2_combout ),
	.Equal131(\router|Equal13~1_combout ),
	.Equal142(\router|Equal14~2_combout ),
	.Equal52(\router|Equal5~2_combout ),
	.Equal91(\router|Equal9~1_combout ),
	.src_channel_0(\router|src_channel[0]~1_combout ),
	.Equal2(\router|Equal2~0_combout ));

spw_babasu_altera_avalon_sc_fifo_18 spill_enable_s1_agent_rdata_fifo(
	.read_latency_shift_reg_0(\spill_enable_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\spill_enable_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_129_0(\spill_enable_s1_agent_rsp_fifo|mem[0][129]~q ),
	.mem_used_01(\spill_enable_s1_agent_rsp_fifo|mem_used[0]~q ),
	.av_readdata_pre_0(\spill_enable_s1_translator|av_readdata_pre[0]~q ),
	.mem_0_0(\spill_enable_s1_agent_rdata_fifo|mem[0][0]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.WideOr0(\rsp_demux_016|WideOr0~0_combout ),
	.clk(clk_clk));

spw_babasu_altera_avalon_sc_fifo_19 spill_enable_s1_agent_rsp_fifo(
	.out_valid_reg(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\spill_enable_s1_agent_rsp_fifo|mem_used[1]~q ),
	.WideOr0(\spill_enable_s1_agent|WideOr0~0_combout ),
	.in_data_reg_68(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ),
	.stateST_UNCOMP_WR_SUBBURST(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.mem_129_0(\spill_enable_s1_agent_rsp_fifo|mem[0][129]~q ),
	.mem_used_0(\spill_enable_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_68_0(\spill_enable_s1_agent_rsp_fifo|mem[0][68]~q ),
	.mem_66_0(\spill_enable_s1_agent_rsp_fifo|mem[0][66]~q ),
	.comb(\spill_enable_s1_agent|comb~0_combout ),
	.mem_130_0(\spill_enable_s1_agent_rsp_fifo|mem[0][130]~q ),
	.mem_78_0(\spill_enable_s1_agent_rsp_fifo|mem[0][78]~q ),
	.mem_77_0(\spill_enable_s1_agent_rsp_fifo|mem[0][77]~q ),
	.mem_76_0(\spill_enable_s1_agent_rsp_fifo|mem[0][76]~q ),
	.mem_75_0(\spill_enable_s1_agent_rsp_fifo|mem[0][75]~q ),
	.mem_74_0(\spill_enable_s1_agent_rsp_fifo|mem[0][74]~q ),
	.mem_105_0(\spill_enable_s1_agent_rsp_fifo|mem[0][105]~q ),
	.mem_106_0(\spill_enable_s1_agent_rsp_fifo|mem[0][106]~q ),
	.mem_107_0(\spill_enable_s1_agent_rsp_fifo|mem[0][107]~q ),
	.mem_108_0(\spill_enable_s1_agent_rsp_fifo|mem[0][108]~q ),
	.mem_109_0(\spill_enable_s1_agent_rsp_fifo|mem[0][109]~q ),
	.mem_110_0(\spill_enable_s1_agent_rsp_fifo|mem[0][110]~q ),
	.mem_111_0(\spill_enable_s1_agent_rsp_fifo|mem[0][111]~q ),
	.mem_112_0(\spill_enable_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_113_0(\spill_enable_s1_agent_rsp_fifo|mem[0][113]~q ),
	.mem_114_0(\spill_enable_s1_agent_rsp_fifo|mem[0][114]~q ),
	.mem_115_0(\spill_enable_s1_agent_rsp_fifo|mem[0][115]~q ),
	.mem_116_0(\spill_enable_s1_agent_rsp_fifo|mem[0][116]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.nxt_out_eop(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.last_packet_beat(\spill_enable_s1_agent|uncompressor|last_packet_beat~2_combout ),
	.WideOr01(\rsp_demux_016|WideOr0~0_combout ),
	.read(\spill_enable_s1_agent_rsp_fifo|read~0_combout ),
	.cp_ready(\spill_enable_s1_agent|cp_ready~3_combout ),
	.in_data_reg_69(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.rf_source_valid(\spill_enable_s1_agent|rf_source_valid~0_combout ),
	.out_byte_cnt_reg_2(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_5(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_4(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_3(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_6(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.sink_ready(\spill_enable_s1_agent|uncompressor|sink_ready~0_combout ),
	.in_data_reg_105(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ),
	.in_data_reg_106(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ),
	.in_data_reg_107(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ),
	.in_data_reg_108(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ),
	.in_data_reg_109(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ),
	.in_data_reg_110(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ),
	.in_data_reg_111(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ),
	.in_data_reg_112(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ),
	.in_data_reg_113(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ),
	.in_data_reg_114(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ),
	.in_data_reg_115(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ),
	.in_data_reg_116(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ),
	.clk(clk_clk));

spw_babasu_altera_avalon_sc_fifo_27 time_out_s1_agent_rsp_fifo(
	.h2f_RREADY_0(h2f_RREADY_0),
	.waitrequest_reset_override(\autostart_s1_translator|waitrequest_reset_override~q ),
	.mem_used_1(\time_out_s1_agent_rsp_fifo|mem_used[1]~q ),
	.in_data_reg_69(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.wait_latency_counter_1(\time_out_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\time_out_s1_translator|wait_latency_counter[0]~q ),
	.nxt_out_eop(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.out_valid_reg(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.stateST_UNCOMP_WR_SUBBURST(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.mem_130_0(\time_out_s1_agent_rsp_fifo|mem[0][130]~q ),
	.empty(\time_out_s1_agent_rdata_fifo|empty~combout ),
	.mem_66_0(\time_out_s1_agent_rsp_fifo|mem[0][66]~q ),
	.mem_used_0(\time_out_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_78_0(\time_out_s1_agent_rsp_fifo|mem[0][78]~q ),
	.mem_77_0(\time_out_s1_agent_rsp_fifo|mem[0][77]~q ),
	.mem_76_0(\time_out_s1_agent_rsp_fifo|mem[0][76]~q ),
	.mem_75_0(\time_out_s1_agent_rsp_fifo|mem[0][75]~q ),
	.mem_74_0(\time_out_s1_agent_rsp_fifo|mem[0][74]~q ),
	.mem_105_0(\time_out_s1_agent_rsp_fifo|mem[0][105]~q ),
	.mem_106_0(\time_out_s1_agent_rsp_fifo|mem[0][106]~q ),
	.mem_107_0(\time_out_s1_agent_rsp_fifo|mem[0][107]~q ),
	.mem_108_0(\time_out_s1_agent_rsp_fifo|mem[0][108]~q ),
	.mem_109_0(\time_out_s1_agent_rsp_fifo|mem[0][109]~q ),
	.mem_110_0(\time_out_s1_agent_rsp_fifo|mem[0][110]~q ),
	.mem_111_0(\time_out_s1_agent_rsp_fifo|mem[0][111]~q ),
	.mem_112_0(\time_out_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_113_0(\time_out_s1_agent_rsp_fifo|mem[0][113]~q ),
	.mem_114_0(\time_out_s1_agent_rsp_fifo|mem[0][114]~q ),
	.mem_115_0(\time_out_s1_agent_rsp_fifo|mem[0][115]~q ),
	.mem_116_0(\time_out_s1_agent_rsp_fifo|mem[0][116]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.last_packet_beat(\time_out_s1_agent|uncompressor|last_packet_beat~2_combout ),
	.write(\time_out_s1_agent_rsp_fifo|write~0_combout ),
	.write1(\time_out_s1_agent_rsp_fifo|write~1_combout ),
	.out_byte_cnt_reg_2(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_6(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.out_uncomp_byte_cnt_reg_5(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_4(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_3(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.in_data_reg_105(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ),
	.in_data_reg_106(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ),
	.in_data_reg_107(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ),
	.in_data_reg_108(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ),
	.in_data_reg_109(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ),
	.in_data_reg_110(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ),
	.in_data_reg_111(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ),
	.in_data_reg_112(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ),
	.in_data_reg_113(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ),
	.in_data_reg_114(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ),
	.in_data_reg_115(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ),
	.in_data_reg_116(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ),
	.clk(clk_clk));

spw_babasu_altera_merlin_slave_agent_13 time_out_s1_agent(
	.h2f_RREADY_0(h2f_RREADY_0),
	.waitrequest_reset_override(\autostart_s1_translator|waitrequest_reset_override~q ),
	.stateST_COMP_TRANS(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.mem_used_1(\time_out_s1_agent_rsp_fifo|mem_used[1]~q ),
	.in_data_reg_69(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.in_narrow_reg(\time_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.wait_latency_counter_1(\time_out_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\time_out_s1_translator|wait_latency_counter[0]~q ),
	.cp_ready(\time_out_s1_agent|cp_ready~0_combout ),
	.cp_ready1(\time_out_s1_agent|cp_ready~1_combout ),
	.empty(\time_out_s1_agent_rdata_fifo|empty~combout ),
	.mem_66_0(\time_out_s1_agent_rsp_fifo|mem[0][66]~q ),
	.mem_used_0(\time_out_s1_agent_rsp_fifo|mem_used[0]~q ),
	.last_packet_beat(\time_out_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.mem_78_0(\time_out_s1_agent_rsp_fifo|mem[0][78]~q ),
	.mem_77_0(\time_out_s1_agent_rsp_fifo|mem[0][77]~q ),
	.mem_76_0(\time_out_s1_agent_rsp_fifo|mem[0][76]~q ),
	.mem_75_0(\time_out_s1_agent_rsp_fifo|mem[0][75]~q ),
	.mem_74_0(\time_out_s1_agent_rsp_fifo|mem[0][74]~q ),
	.last_packet_beat1(\time_out_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.last_packet_beat2(\time_out_s1_agent|uncompressor|last_packet_beat~2_combout ),
	.cp_ready2(\time_out_s1_agent|cp_ready~2_combout ),
	.clk_clk(clk_clk));

spw_babasu_altera_avalon_sc_fifo_22 tick_out_s1_agent_rdata_fifo(
	.h2f_RREADY_0(h2f_RREADY_0),
	.read_latency_shift_reg_0(\tick_out_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\tick_out_s1_agent_rdata_fifo|mem_used[0]~q ),
	.empty1(\tick_out_s1_agent_rdata_fifo|empty~combout ),
	.av_readdata_pre_0(\tick_out_s1_translator|av_readdata_pre[0]~q ),
	.mem_0_0(\tick_out_s1_agent_rdata_fifo|mem[0][0]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.clk(clk_clk));

spw_babasu_altera_avalon_sc_fifo_23 tick_out_s1_agent_rsp_fifo(
	.h2f_RREADY_0(h2f_RREADY_0),
	.waitrequest_reset_override(\autostart_s1_translator|waitrequest_reset_override~q ),
	.mem_used_1(\tick_out_s1_agent_rsp_fifo|mem_used[1]~q ),
	.in_data_reg_69(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.wait_latency_counter_1(\tick_out_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\tick_out_s1_translator|wait_latency_counter[0]~q ),
	.nxt_out_eop(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.out_valid_reg(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.stateST_UNCOMP_WR_SUBBURST(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.mem_130_0(\tick_out_s1_agent_rsp_fifo|mem[0][130]~q ),
	.empty(\tick_out_s1_agent_rdata_fifo|empty~combout ),
	.mem_66_0(\tick_out_s1_agent_rsp_fifo|mem[0][66]~q ),
	.mem_used_0(\tick_out_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_78_0(\tick_out_s1_agent_rsp_fifo|mem[0][78]~q ),
	.mem_77_0(\tick_out_s1_agent_rsp_fifo|mem[0][77]~q ),
	.mem_76_0(\tick_out_s1_agent_rsp_fifo|mem[0][76]~q ),
	.mem_75_0(\tick_out_s1_agent_rsp_fifo|mem[0][75]~q ),
	.mem_74_0(\tick_out_s1_agent_rsp_fifo|mem[0][74]~q ),
	.mem_105_0(\tick_out_s1_agent_rsp_fifo|mem[0][105]~q ),
	.mem_106_0(\tick_out_s1_agent_rsp_fifo|mem[0][106]~q ),
	.mem_107_0(\tick_out_s1_agent_rsp_fifo|mem[0][107]~q ),
	.mem_108_0(\tick_out_s1_agent_rsp_fifo|mem[0][108]~q ),
	.mem_109_0(\tick_out_s1_agent_rsp_fifo|mem[0][109]~q ),
	.mem_110_0(\tick_out_s1_agent_rsp_fifo|mem[0][110]~q ),
	.mem_111_0(\tick_out_s1_agent_rsp_fifo|mem[0][111]~q ),
	.mem_112_0(\tick_out_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_113_0(\tick_out_s1_agent_rsp_fifo|mem[0][113]~q ),
	.mem_114_0(\tick_out_s1_agent_rsp_fifo|mem[0][114]~q ),
	.mem_115_0(\tick_out_s1_agent_rsp_fifo|mem[0][115]~q ),
	.mem_116_0(\tick_out_s1_agent_rsp_fifo|mem[0][116]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.last_packet_beat(\tick_out_s1_agent|uncompressor|last_packet_beat~2_combout ),
	.write(\tick_out_s1_agent_rsp_fifo|write~0_combout ),
	.write1(\tick_out_s1_agent_rsp_fifo|write~1_combout ),
	.out_byte_cnt_reg_2(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_3(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_4(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_5(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_6(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.in_data_reg_105(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ),
	.in_data_reg_106(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ),
	.in_data_reg_107(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ),
	.in_data_reg_108(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ),
	.in_data_reg_109(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ),
	.in_data_reg_110(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ),
	.in_data_reg_111(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ),
	.in_data_reg_112(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ),
	.in_data_reg_113(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ),
	.in_data_reg_114(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ),
	.in_data_reg_115(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ),
	.in_data_reg_116(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ),
	.clk(clk_clk));

spw_babasu_altera_merlin_slave_agent_11 tick_out_s1_agent(
	.h2f_RREADY_0(h2f_RREADY_0),
	.waitrequest_reset_override(\autostart_s1_translator|waitrequest_reset_override~q ),
	.stateST_COMP_TRANS(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.mem_used_1(\tick_out_s1_agent_rsp_fifo|mem_used[1]~q ),
	.in_data_reg_69(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.in_narrow_reg(\tick_out_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.wait_latency_counter_1(\tick_out_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\tick_out_s1_translator|wait_latency_counter[0]~q ),
	.cp_ready(\tick_out_s1_agent|cp_ready~0_combout ),
	.cp_ready1(\tick_out_s1_agent|cp_ready~1_combout ),
	.empty(\tick_out_s1_agent_rdata_fifo|empty~combout ),
	.mem_66_0(\tick_out_s1_agent_rsp_fifo|mem[0][66]~q ),
	.mem_used_0(\tick_out_s1_agent_rsp_fifo|mem_used[0]~q ),
	.last_packet_beat(\tick_out_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.mem_78_0(\tick_out_s1_agent_rsp_fifo|mem[0][78]~q ),
	.mem_77_0(\tick_out_s1_agent_rsp_fifo|mem[0][77]~q ),
	.mem_76_0(\tick_out_s1_agent_rsp_fifo|mem[0][76]~q ),
	.mem_75_0(\tick_out_s1_agent_rsp_fifo|mem[0][75]~q ),
	.mem_74_0(\tick_out_s1_agent_rsp_fifo|mem[0][74]~q ),
	.last_packet_beat1(\tick_out_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.last_packet_beat2(\tick_out_s1_agent|uncompressor|last_packet_beat~2_combout ),
	.cp_ready2(\tick_out_s1_agent|cp_ready~2_combout ),
	.clk_clk(clk_clk));

spw_babasu_altera_avalon_sc_fifo_16 rx_empty_s1_agent_rdata_fifo(
	.h2f_RREADY_0(h2f_RREADY_0),
	.read_latency_shift_reg_0(\rx_empty_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\rx_empty_s1_agent_rdata_fifo|mem_used[0]~q ),
	.empty1(\rx_empty_s1_agent_rdata_fifo|empty~combout ),
	.av_readdata_pre_0(\rx_empty_s1_translator|av_readdata_pre[0]~q ),
	.mem_0_0(\rx_empty_s1_agent_rdata_fifo|mem[0][0]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.clk(clk_clk));

spw_babasu_altera_merlin_slave_agent_2 data_i_s1_agent(
	.waitrequest_reset_override(\autostart_s1_translator|waitrequest_reset_override~q ),
	.stateST_COMP_TRANS(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.out_valid_reg(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\data_i_s1_agent_rsp_fifo|mem_used[1]~q ),
	.in_narrow_reg(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.in_byteen_reg_3(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ),
	.in_byteen_reg_2(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ),
	.in_byteen_reg_1(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ),
	.in_byteen_reg_0(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ),
	.WideOr0(\data_i_s1_agent|WideOr0~0_combout ),
	.wait_latency_counter_1(wait_latency_counter_15),
	.wait_latency_counter_0(wait_latency_counter_05),
	.in_data_reg_68(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ),
	.cp_ready(\data_i_s1_agent|cp_ready~0_combout ),
	.read_latency_shift_reg_0(\data_i_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\data_i_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_129_0(\data_i_s1_agent_rsp_fifo|mem[0][129]~q ),
	.mem_used_01(\data_i_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_66_0(\data_i_s1_agent_rsp_fifo|mem[0][66]~q ),
	.comb(\data_i_s1_agent|comb~0_combout ),
	.last_packet_beat(\data_i_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.mem_78_0(\data_i_s1_agent_rsp_fifo|mem[0][78]~q ),
	.mem_77_0(\data_i_s1_agent_rsp_fifo|mem[0][77]~q ),
	.mem_76_0(\data_i_s1_agent_rsp_fifo|mem[0][76]~q ),
	.mem_75_0(\data_i_s1_agent_rsp_fifo|mem[0][75]~q ),
	.mem_74_0(\data_i_s1_agent_rsp_fifo|mem[0][74]~q ),
	.last_packet_beat1(\data_i_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.m0_write1(m0_write1),
	.nxt_out_eop(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.cp_ready1(\data_i_s1_agent|cp_ready~3_combout ),
	.last_packet_beat2(\data_i_s1_agent|uncompressor|last_packet_beat~2_combout ),
	.WideOr01(\rsp_demux_005|WideOr0~0_combout ),
	.read(\data_i_s1_agent_rsp_fifo|read~0_combout ),
	.cp_ready2(\data_i_s1_agent|cp_ready~4_combout ),
	.in_data_reg_69(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.rf_source_valid(\data_i_s1_agent|rf_source_valid~0_combout ),
	.rf_sink_ready(\data_i_s1_agent|uncompressor|sink_ready~0_combout ),
	.clk_clk(clk_clk));

spw_babasu_altera_avalon_sc_fifo_8 flags_s1_agent_rdata_fifo(
	.h2f_RREADY_0(h2f_RREADY_0),
	.read_latency_shift_reg_0(\flags_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\flags_s1_agent_rdata_fifo|mem_used[0]~q ),
	.empty1(\flags_s1_agent_rdata_fifo|empty~combout ),
	.av_readdata_pre_0(\flags_s1_translator|av_readdata_pre[0]~q ),
	.mem_0_0(\flags_s1_agent_rdata_fifo|mem[0][0]~q ),
	.mem_1_0(\flags_s1_agent_rdata_fifo|mem[0][1]~q ),
	.av_readdata_pre_1(\flags_s1_translator|av_readdata_pre[1]~q ),
	.mem_2_0(\flags_s1_agent_rdata_fifo|mem[0][2]~q ),
	.av_readdata_pre_2(\flags_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\flags_s1_translator|av_readdata_pre[3]~q ),
	.mem_3_0(\flags_s1_agent_rdata_fifo|mem[0][3]~q ),
	.av_readdata_pre_4(\flags_s1_translator|av_readdata_pre[4]~q ),
	.mem_4_0(\flags_s1_agent_rdata_fifo|mem[0][4]~q ),
	.av_readdata_pre_5(\flags_s1_translator|av_readdata_pre[5]~q ),
	.mem_5_0(\flags_s1_agent_rdata_fifo|mem[0][5]~q ),
	.av_readdata_pre_6(\flags_s1_translator|av_readdata_pre[6]~q ),
	.mem_6_0(\flags_s1_agent_rdata_fifo|mem[0][6]~q ),
	.av_readdata_pre_7(\flags_s1_translator|av_readdata_pre[7]~q ),
	.mem_7_0(\flags_s1_agent_rdata_fifo|mem[0][7]~q ),
	.mem_8_0(\flags_s1_agent_rdata_fifo|mem[0][8]~q ),
	.av_readdata_pre_8(\flags_s1_translator|av_readdata_pre[8]~q ),
	.mem_9_0(\flags_s1_agent_rdata_fifo|mem[0][9]~q ),
	.av_readdata_pre_9(\flags_s1_translator|av_readdata_pre[9]~q ),
	.mem_10_0(\flags_s1_agent_rdata_fifo|mem[0][10]~q ),
	.av_readdata_pre_10(\flags_s1_translator|av_readdata_pre[10]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.clk(clk_clk));

spw_babasu_altera_avalon_sc_fifo_9 flags_s1_agent_rsp_fifo(
	.h2f_RREADY_0(h2f_RREADY_0),
	.waitrequest_reset_override(\autostart_s1_translator|waitrequest_reset_override~q ),
	.in_data_reg_69(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.mem_used_1(\flags_s1_agent_rsp_fifo|mem_used[1]~q ),
	.wait_latency_counter_1(\flags_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\flags_s1_translator|wait_latency_counter[0]~q ),
	.out_valid_reg(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.stateST_UNCOMP_WR_SUBBURST(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.empty(\flags_s1_agent_rdata_fifo|empty~combout ),
	.mem_66_0(\flags_s1_agent_rsp_fifo|mem[0][66]~q ),
	.mem_used_0(\flags_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_78_0(\flags_s1_agent_rsp_fifo|mem[0][78]~q ),
	.mem_77_0(\flags_s1_agent_rsp_fifo|mem[0][77]~q ),
	.mem_76_0(\flags_s1_agent_rsp_fifo|mem[0][76]~q ),
	.mem_75_0(\flags_s1_agent_rsp_fifo|mem[0][75]~q ),
	.mem_74_0(\flags_s1_agent_rsp_fifo|mem[0][74]~q ),
	.last_packet_beat(\flags_s1_agent|uncompressor|last_packet_beat~3_combout ),
	.mem_130_0(\flags_s1_agent_rsp_fifo|mem[0][130]~q ),
	.mem_105_0(\flags_s1_agent_rsp_fifo|mem[0][105]~q ),
	.mem_106_0(\flags_s1_agent_rsp_fifo|mem[0][106]~q ),
	.mem_107_0(\flags_s1_agent_rsp_fifo|mem[0][107]~q ),
	.mem_108_0(\flags_s1_agent_rsp_fifo|mem[0][108]~q ),
	.mem_109_0(\flags_s1_agent_rsp_fifo|mem[0][109]~q ),
	.mem_110_0(\flags_s1_agent_rsp_fifo|mem[0][110]~q ),
	.mem_111_0(\flags_s1_agent_rsp_fifo|mem[0][111]~q ),
	.mem_112_0(\flags_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_113_0(\flags_s1_agent_rsp_fifo|mem[0][113]~q ),
	.mem_114_0(\flags_s1_agent_rsp_fifo|mem[0][114]~q ),
	.mem_115_0(\flags_s1_agent_rsp_fifo|mem[0][115]~q ),
	.mem_116_0(\flags_s1_agent_rsp_fifo|mem[0][116]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.nxt_out_eop(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.out_byte_cnt_reg_2(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.write(\flags_s1_agent_rsp_fifo|write~0_combout ),
	.write1(\flags_s1_agent_rsp_fifo|write~1_combout ),
	.out_uncomp_byte_cnt_reg_6(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.out_uncomp_byte_cnt_reg_5(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_4(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_3(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.in_data_reg_105(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ),
	.in_data_reg_106(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ),
	.in_data_reg_107(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ),
	.in_data_reg_108(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ),
	.in_data_reg_109(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ),
	.in_data_reg_110(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ),
	.in_data_reg_111(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ),
	.in_data_reg_112(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ),
	.in_data_reg_113(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ),
	.in_data_reg_114(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ),
	.in_data_reg_115(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ),
	.in_data_reg_116(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ),
	.clk(clk_clk));

spw_babasu_altera_merlin_slave_agent_4 flags_s1_agent(
	.h2f_RREADY_0(h2f_RREADY_0),
	.waitrequest_reset_override(\autostart_s1_translator|waitrequest_reset_override~q ),
	.in_data_reg_69(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.stateST_COMP_TRANS(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.in_narrow_reg(\flags_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.wait_latency_counter_1(\flags_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\flags_s1_translator|wait_latency_counter[0]~q ),
	.cp_ready(\flags_s1_agent|cp_ready~0_combout ),
	.empty(\flags_s1_agent_rdata_fifo|empty~combout ),
	.mem_66_0(\flags_s1_agent_rsp_fifo|mem[0][66]~q ),
	.mem_used_0(\flags_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_78_0(\flags_s1_agent_rsp_fifo|mem[0][78]~q ),
	.mem_77_0(\flags_s1_agent_rsp_fifo|mem[0][77]~q ),
	.mem_76_0(\flags_s1_agent_rsp_fifo|mem[0][76]~q ),
	.mem_75_0(\flags_s1_agent_rsp_fifo|mem[0][75]~q ),
	.mem_74_0(\flags_s1_agent_rsp_fifo|mem[0][74]~q ),
	.last_packet_beat(\flags_s1_agent|uncompressor|last_packet_beat~3_combout ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.cp_ready1(\flags_s1_agent|cp_ready~1_combout ),
	.clk_clk(clk_clk));

spw_babasu_altera_avalon_sc_fifo_2 currentstate_s1_agent_rdata_fifo(
	.h2f_RREADY_0(h2f_RREADY_0),
	.read_latency_shift_reg_0(\currentstate_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\currentstate_s1_agent_rdata_fifo|mem_used[0]~q ),
	.empty1(\currentstate_s1_agent_rdata_fifo|empty~combout ),
	.av_readdata_pre_0(\currentstate_s1_translator|av_readdata_pre[0]~q ),
	.mem_0_0(\currentstate_s1_agent_rdata_fifo|mem[0][0]~q ),
	.av_readdata_pre_1(\currentstate_s1_translator|av_readdata_pre[1]~q ),
	.mem_1_0(\currentstate_s1_agent_rdata_fifo|mem[0][1]~q ),
	.av_readdata_pre_2(\currentstate_s1_translator|av_readdata_pre[2]~q ),
	.mem_2_0(\currentstate_s1_agent_rdata_fifo|mem[0][2]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.clk(clk_clk));

spw_babasu_altera_avalon_sc_fifo_3 currentstate_s1_agent_rsp_fifo(
	.h2f_RREADY_0(h2f_RREADY_0),
	.waitrequest_reset_override(\autostart_s1_translator|waitrequest_reset_override~q ),
	.mem_used_1(\currentstate_s1_agent_rsp_fifo|mem_used[1]~q ),
	.in_data_reg_69(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.wait_latency_counter_1(\currentstate_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\currentstate_s1_translator|wait_latency_counter[0]~q ),
	.nxt_out_eop(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.out_valid_reg(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.stateST_UNCOMP_WR_SUBBURST(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.mem_130_0(\currentstate_s1_agent_rsp_fifo|mem[0][130]~q ),
	.empty(\currentstate_s1_agent_rdata_fifo|empty~combout ),
	.mem_66_0(\currentstate_s1_agent_rsp_fifo|mem[0][66]~q ),
	.mem_used_0(\currentstate_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_78_0(\currentstate_s1_agent_rsp_fifo|mem[0][78]~q ),
	.mem_77_0(\currentstate_s1_agent_rsp_fifo|mem[0][77]~q ),
	.mem_76_0(\currentstate_s1_agent_rsp_fifo|mem[0][76]~q ),
	.mem_75_0(\currentstate_s1_agent_rsp_fifo|mem[0][75]~q ),
	.mem_74_0(\currentstate_s1_agent_rsp_fifo|mem[0][74]~q ),
	.mem_105_0(\currentstate_s1_agent_rsp_fifo|mem[0][105]~q ),
	.mem_106_0(\currentstate_s1_agent_rsp_fifo|mem[0][106]~q ),
	.mem_107_0(\currentstate_s1_agent_rsp_fifo|mem[0][107]~q ),
	.mem_108_0(\currentstate_s1_agent_rsp_fifo|mem[0][108]~q ),
	.mem_109_0(\currentstate_s1_agent_rsp_fifo|mem[0][109]~q ),
	.mem_110_0(\currentstate_s1_agent_rsp_fifo|mem[0][110]~q ),
	.mem_111_0(\currentstate_s1_agent_rsp_fifo|mem[0][111]~q ),
	.mem_112_0(\currentstate_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_113_0(\currentstate_s1_agent_rsp_fifo|mem[0][113]~q ),
	.mem_114_0(\currentstate_s1_agent_rsp_fifo|mem[0][114]~q ),
	.mem_115_0(\currentstate_s1_agent_rsp_fifo|mem[0][115]~q ),
	.mem_116_0(\currentstate_s1_agent_rsp_fifo|mem[0][116]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.last_packet_beat(\currentstate_s1_agent|uncompressor|last_packet_beat~2_combout ),
	.write(\currentstate_s1_agent_rsp_fifo|write~0_combout ),
	.write1(\currentstate_s1_agent_rsp_fifo|write~1_combout ),
	.out_byte_cnt_reg_2(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_3(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_4(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_5(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_6(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.in_data_reg_105(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ),
	.in_data_reg_106(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ),
	.in_data_reg_107(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ),
	.in_data_reg_108(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ),
	.in_data_reg_109(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ),
	.in_data_reg_110(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ),
	.in_data_reg_111(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ),
	.in_data_reg_112(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ),
	.in_data_reg_113(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ),
	.in_data_reg_114(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ),
	.in_data_reg_115(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ),
	.in_data_reg_116(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ),
	.clk(clk_clk));

spw_babasu_altera_merlin_slave_agent_1 currentstate_s1_agent(
	.h2f_RREADY_0(h2f_RREADY_0),
	.waitrequest_reset_override(\autostart_s1_translator|waitrequest_reset_override~q ),
	.stateST_COMP_TRANS(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.mem_used_1(\currentstate_s1_agent_rsp_fifo|mem_used[1]~q ),
	.in_data_reg_69(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.in_narrow_reg(\currentstate_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.wait_latency_counter_1(\currentstate_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\currentstate_s1_translator|wait_latency_counter[0]~q ),
	.cp_ready(\currentstate_s1_agent|cp_ready~0_combout ),
	.cp_ready1(\currentstate_s1_agent|cp_ready~1_combout ),
	.empty(\currentstate_s1_agent_rdata_fifo|empty~combout ),
	.mem_66_0(\currentstate_s1_agent_rsp_fifo|mem[0][66]~q ),
	.mem_used_0(\currentstate_s1_agent_rsp_fifo|mem_used[0]~q ),
	.last_packet_beat(\currentstate_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.mem_78_0(\currentstate_s1_agent_rsp_fifo|mem[0][78]~q ),
	.mem_77_0(\currentstate_s1_agent_rsp_fifo|mem[0][77]~q ),
	.mem_76_0(\currentstate_s1_agent_rsp_fifo|mem[0][76]~q ),
	.mem_75_0(\currentstate_s1_agent_rsp_fifo|mem[0][75]~q ),
	.mem_74_0(\currentstate_s1_agent_rsp_fifo|mem[0][74]~q ),
	.last_packet_beat1(\currentstate_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.last_packet_beat2(\currentstate_s1_agent|uncompressor|last_packet_beat~2_combout ),
	.cp_ready2(\currentstate_s1_agent|cp_ready~2_combout ),
	.clk_clk(clk_clk));

spw_babasu_altera_avalon_sc_fifo autostart_s1_agent_rdata_fifo(
	.read_latency_shift_reg_0(\autostart_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\autostart_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_129_0(\autostart_s1_agent_rsp_fifo|mem[0][129]~q ),
	.mem_used_01(\autostart_s1_agent_rsp_fifo|mem_used[0]~q ),
	.av_readdata_pre_0(\autostart_s1_translator|av_readdata_pre[0]~q ),
	.mem_0_0(\autostart_s1_agent_rdata_fifo|mem[0][0]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.WideOr0(\rsp_demux_002|WideOr0~0_combout ),
	.clk(clk_clk));

spw_babasu_altera_avalon_sc_fifo_1 autostart_s1_agent_rsp_fifo(
	.out_valid_reg(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\autostart_s1_agent_rsp_fifo|mem_used[1]~q ),
	.WideOr0(\autostart_s1_agent|WideOr0~0_combout ),
	.in_data_reg_68(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ),
	.stateST_UNCOMP_WR_SUBBURST(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.mem_129_0(\autostart_s1_agent_rsp_fifo|mem[0][129]~q ),
	.mem_used_0(\autostart_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_68_0(\autostart_s1_agent_rsp_fifo|mem[0][68]~q ),
	.mem_66_0(\autostart_s1_agent_rsp_fifo|mem[0][66]~q ),
	.comb(\autostart_s1_agent|comb~0_combout ),
	.mem_130_0(\autostart_s1_agent_rsp_fifo|mem[0][130]~q ),
	.mem_78_0(\autostart_s1_agent_rsp_fifo|mem[0][78]~q ),
	.mem_77_0(\autostart_s1_agent_rsp_fifo|mem[0][77]~q ),
	.mem_76_0(\autostart_s1_agent_rsp_fifo|mem[0][76]~q ),
	.mem_75_0(\autostart_s1_agent_rsp_fifo|mem[0][75]~q ),
	.mem_74_0(\autostart_s1_agent_rsp_fifo|mem[0][74]~q ),
	.mem_105_0(\autostart_s1_agent_rsp_fifo|mem[0][105]~q ),
	.mem_106_0(\autostart_s1_agent_rsp_fifo|mem[0][106]~q ),
	.mem_107_0(\autostart_s1_agent_rsp_fifo|mem[0][107]~q ),
	.mem_108_0(\autostart_s1_agent_rsp_fifo|mem[0][108]~q ),
	.mem_109_0(\autostart_s1_agent_rsp_fifo|mem[0][109]~q ),
	.mem_110_0(\autostart_s1_agent_rsp_fifo|mem[0][110]~q ),
	.mem_111_0(\autostart_s1_agent_rsp_fifo|mem[0][111]~q ),
	.mem_112_0(\autostart_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_113_0(\autostart_s1_agent_rsp_fifo|mem[0][113]~q ),
	.mem_114_0(\autostart_s1_agent_rsp_fifo|mem[0][114]~q ),
	.mem_115_0(\autostart_s1_agent_rsp_fifo|mem[0][115]~q ),
	.mem_116_0(\autostart_s1_agent_rsp_fifo|mem[0][116]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.nxt_out_eop(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.last_packet_beat(\autostart_s1_agent|uncompressor|last_packet_beat~2_combout ),
	.WideOr01(\rsp_demux_002|WideOr0~0_combout ),
	.read(\autostart_s1_agent_rsp_fifo|read~0_combout ),
	.cp_ready(\autostart_s1_agent|cp_ready~4_combout ),
	.in_data_reg_69(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.rf_source_valid(\autostart_s1_agent|rf_source_valid~0_combout ),
	.out_byte_cnt_reg_2(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_5(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_4(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_3(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_6(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.sink_ready(\autostart_s1_agent|uncompressor|sink_ready~0_combout ),
	.in_data_reg_105(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ),
	.in_data_reg_106(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ),
	.in_data_reg_107(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ),
	.in_data_reg_108(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ),
	.in_data_reg_109(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ),
	.in_data_reg_110(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ),
	.in_data_reg_111(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ),
	.in_data_reg_112(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ),
	.in_data_reg_113(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ),
	.in_data_reg_114(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ),
	.in_data_reg_115(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ),
	.in_data_reg_116(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ),
	.clk(clk_clk));

spw_babasu_altera_merlin_slave_agent autostart_s1_agent(
	.waitrequest_reset_override(\autostart_s1_translator|waitrequest_reset_override~q ),
	.stateST_COMP_TRANS(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.out_valid_reg(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\autostart_s1_agent_rsp_fifo|mem_used[1]~q ),
	.in_narrow_reg(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.in_byteen_reg_3(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ),
	.in_byteen_reg_2(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ),
	.in_byteen_reg_1(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ),
	.in_byteen_reg_0(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ),
	.WideOr0(\autostart_s1_agent|WideOr0~0_combout ),
	.wait_latency_counter_1(wait_latency_counter_18),
	.wait_latency_counter_0(wait_latency_counter_08),
	.in_data_reg_68(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ),
	.cp_ready(\autostart_s1_agent|cp_ready~0_combout ),
	.read_latency_shift_reg_0(\autostart_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\autostart_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_129_0(\autostart_s1_agent_rsp_fifo|mem[0][129]~q ),
	.mem_used_01(\autostart_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_66_0(\autostart_s1_agent_rsp_fifo|mem[0][66]~q ),
	.comb(\autostart_s1_agent|comb~0_combout ),
	.last_packet_beat(\autostart_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.mem_78_0(\autostart_s1_agent_rsp_fifo|mem[0][78]~q ),
	.mem_77_0(\autostart_s1_agent_rsp_fifo|mem[0][77]~q ),
	.mem_76_0(\autostart_s1_agent_rsp_fifo|mem[0][76]~q ),
	.mem_75_0(\autostart_s1_agent_rsp_fifo|mem[0][75]~q ),
	.mem_74_0(\autostart_s1_agent_rsp_fifo|mem[0][74]~q ),
	.last_packet_beat1(\autostart_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.m0_write1(m0_write),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.nxt_out_eop(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.cp_ready1(\autostart_s1_agent|cp_ready~3_combout ),
	.last_packet_beat2(\autostart_s1_agent|uncompressor|last_packet_beat~2_combout ),
	.WideOr01(\rsp_demux_002|WideOr0~0_combout ),
	.read(\autostart_s1_agent_rsp_fifo|read~0_combout ),
	.cp_ready2(\autostart_s1_agent|cp_ready~4_combout ),
	.in_data_reg_69(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.rf_source_valid(\autostart_s1_agent|rf_source_valid~0_combout ),
	.rf_sink_ready(\autostart_s1_agent|uncompressor|sink_ready~0_combout ),
	.clk_clk(clk_clk));

spw_babasu_altera_avalon_sc_fifo_10 link_disable_s1_agent_rdata_fifo(
	.read_latency_shift_reg_0(\link_disable_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\link_disable_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_129_0(\link_disable_s1_agent_rsp_fifo|mem[0][129]~q ),
	.mem_used_01(\link_disable_s1_agent_rsp_fifo|mem_used[0]~q ),
	.av_readdata_pre_0(\link_disable_s1_translator|av_readdata_pre[0]~q ),
	.mem_0_0(\link_disable_s1_agent_rdata_fifo|mem[0][0]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.WideOr0(\rsp_demux_001|WideOr0~0_combout ),
	.clk(clk_clk));

spw_babasu_altera_merlin_slave_agent_15 tx_full_s1_agent(
	.h2f_RREADY_0(h2f_RREADY_0),
	.waitrequest_reset_override(\autostart_s1_translator|waitrequest_reset_override~q ),
	.in_data_reg_69(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.stateST_COMP_TRANS(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.in_narrow_reg(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.wait_latency_counter_1(\tx_full_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\tx_full_s1_translator|wait_latency_counter[0]~q ),
	.cp_ready(\tx_full_s1_agent|cp_ready~0_combout ),
	.empty(\tx_full_s1_agent_rdata_fifo|empty~combout ),
	.mem_66_0(\tx_full_s1_agent_rsp_fifo|mem[0][66]~q ),
	.mem_used_0(\tx_full_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_78_0(\tx_full_s1_agent_rsp_fifo|mem[0][78]~q ),
	.mem_77_0(\tx_full_s1_agent_rsp_fifo|mem[0][77]~q ),
	.mem_76_0(\tx_full_s1_agent_rsp_fifo|mem[0][76]~q ),
	.mem_75_0(\tx_full_s1_agent_rsp_fifo|mem[0][75]~q ),
	.mem_74_0(\tx_full_s1_agent_rsp_fifo|mem[0][74]~q ),
	.last_packet_beat(\tx_full_s1_agent|uncompressor|last_packet_beat~3_combout ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.cp_ready1(\tx_full_s1_agent|cp_ready~1_combout ),
	.clk_clk(clk_clk));

spw_babasu_altera_avalon_sc_fifo_32 wr_data_s1_agent_rdata_fifo(
	.read_latency_shift_reg_0(\wr_data_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\wr_data_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_129_0(\wr_data_s1_agent_rsp_fifo|mem[0][129]~q ),
	.mem_used_01(\wr_data_s1_agent_rsp_fifo|mem_used[0]~q ),
	.av_readdata_pre_0(\wr_data_s1_translator|av_readdata_pre[0]~q ),
	.mem_0_0(\wr_data_s1_agent_rdata_fifo|mem[0][0]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.WideOr0(\rsp_demux_006|WideOr0~0_combout ),
	.clk(clk_clk));

spw_babasu_altera_avalon_sc_fifo_33 wr_data_s1_agent_rsp_fifo(
	.out_valid_reg(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\wr_data_s1_agent_rsp_fifo|mem_used[1]~q ),
	.WideOr0(\wr_data_s1_agent|WideOr0~0_combout ),
	.in_data_reg_68(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ),
	.stateST_UNCOMP_WR_SUBBURST(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.mem_129_0(\wr_data_s1_agent_rsp_fifo|mem[0][129]~q ),
	.mem_used_0(\wr_data_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_68_0(\wr_data_s1_agent_rsp_fifo|mem[0][68]~q ),
	.mem_66_0(\wr_data_s1_agent_rsp_fifo|mem[0][66]~q ),
	.comb(\wr_data_s1_agent|comb~0_combout ),
	.mem_130_0(\wr_data_s1_agent_rsp_fifo|mem[0][130]~q ),
	.mem_78_0(\wr_data_s1_agent_rsp_fifo|mem[0][78]~q ),
	.mem_77_0(\wr_data_s1_agent_rsp_fifo|mem[0][77]~q ),
	.mem_76_0(\wr_data_s1_agent_rsp_fifo|mem[0][76]~q ),
	.mem_75_0(\wr_data_s1_agent_rsp_fifo|mem[0][75]~q ),
	.mem_74_0(\wr_data_s1_agent_rsp_fifo|mem[0][74]~q ),
	.mem_105_0(\wr_data_s1_agent_rsp_fifo|mem[0][105]~q ),
	.mem_106_0(\wr_data_s1_agent_rsp_fifo|mem[0][106]~q ),
	.mem_107_0(\wr_data_s1_agent_rsp_fifo|mem[0][107]~q ),
	.mem_108_0(\wr_data_s1_agent_rsp_fifo|mem[0][108]~q ),
	.mem_109_0(\wr_data_s1_agent_rsp_fifo|mem[0][109]~q ),
	.mem_110_0(\wr_data_s1_agent_rsp_fifo|mem[0][110]~q ),
	.mem_111_0(\wr_data_s1_agent_rsp_fifo|mem[0][111]~q ),
	.mem_112_0(\wr_data_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_113_0(\wr_data_s1_agent_rsp_fifo|mem[0][113]~q ),
	.mem_114_0(\wr_data_s1_agent_rsp_fifo|mem[0][114]~q ),
	.mem_115_0(\wr_data_s1_agent_rsp_fifo|mem[0][115]~q ),
	.mem_116_0(\wr_data_s1_agent_rsp_fifo|mem[0][116]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.nxt_out_eop(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.last_packet_beat(\wr_data_s1_agent|uncompressor|last_packet_beat~2_combout ),
	.WideOr01(\rsp_demux_006|WideOr0~0_combout ),
	.read(\wr_data_s1_agent_rsp_fifo|read~0_combout ),
	.cp_ready(\wr_data_s1_agent|cp_ready~4_combout ),
	.in_data_reg_69(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.rf_source_valid(\wr_data_s1_agent|rf_source_valid~0_combout ),
	.out_byte_cnt_reg_2(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_4(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_3(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_5(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_6(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.sink_ready(\wr_data_s1_agent|uncompressor|sink_ready~0_combout ),
	.in_data_reg_105(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ),
	.in_data_reg_106(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ),
	.in_data_reg_107(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ),
	.in_data_reg_108(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ),
	.in_data_reg_109(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ),
	.in_data_reg_110(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ),
	.in_data_reg_111(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ),
	.in_data_reg_112(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ),
	.in_data_reg_113(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ),
	.in_data_reg_114(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ),
	.in_data_reg_115(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ),
	.in_data_reg_116(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ),
	.clk(clk_clk));

spw_babasu_altera_merlin_slave_agent_16 wr_data_s1_agent(
	.waitrequest_reset_override(\autostart_s1_translator|waitrequest_reset_override~q ),
	.stateST_COMP_TRANS(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.out_valid_reg(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\wr_data_s1_agent_rsp_fifo|mem_used[1]~q ),
	.in_narrow_reg(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.in_byteen_reg_3(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ),
	.in_byteen_reg_2(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ),
	.in_byteen_reg_1(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ),
	.in_byteen_reg_0(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ),
	.WideOr0(\wr_data_s1_agent|WideOr0~0_combout ),
	.wait_latency_counter_1(wait_latency_counter_19),
	.wait_latency_counter_0(wait_latency_counter_09),
	.in_data_reg_68(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ),
	.cp_ready(\wr_data_s1_agent|cp_ready~0_combout ),
	.read_latency_shift_reg_0(\wr_data_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\wr_data_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_129_0(\wr_data_s1_agent_rsp_fifo|mem[0][129]~q ),
	.mem_used_01(\wr_data_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_66_0(\wr_data_s1_agent_rsp_fifo|mem[0][66]~q ),
	.comb(\wr_data_s1_agent|comb~0_combout ),
	.last_packet_beat(\wr_data_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.mem_78_0(\wr_data_s1_agent_rsp_fifo|mem[0][78]~q ),
	.mem_77_0(\wr_data_s1_agent_rsp_fifo|mem[0][77]~q ),
	.mem_76_0(\wr_data_s1_agent_rsp_fifo|mem[0][76]~q ),
	.mem_75_0(\wr_data_s1_agent_rsp_fifo|mem[0][75]~q ),
	.mem_74_0(\wr_data_s1_agent_rsp_fifo|mem[0][74]~q ),
	.last_packet_beat1(\wr_data_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.m0_write1(m0_write9),
	.nxt_out_eop(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.cp_ready1(\wr_data_s1_agent|cp_ready~3_combout ),
	.last_packet_beat2(\wr_data_s1_agent|uncompressor|last_packet_beat~2_combout ),
	.WideOr01(\rsp_demux_006|WideOr0~0_combout ),
	.read(\wr_data_s1_agent_rsp_fifo|read~0_combout ),
	.cp_ready2(\wr_data_s1_agent|cp_ready~4_combout ),
	.in_data_reg_69(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.rf_source_valid(\wr_data_s1_agent|rf_source_valid~0_combout ),
	.rf_sink_ready(\wr_data_s1_agent|uncompressor|sink_ready~0_combout ),
	.clk_clk(clk_clk));

spw_babasu_altera_avalon_sc_fifo_4 data_i_s1_agent_rdata_fifo(
	.read_latency_shift_reg_0(\data_i_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\data_i_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_129_0(\data_i_s1_agent_rsp_fifo|mem[0][129]~q ),
	.mem_used_01(\data_i_s1_agent_rsp_fifo|mem_used[0]~q ),
	.av_readdata_pre_0(\data_i_s1_translator|av_readdata_pre[0]~q ),
	.always4(\data_i_s1_agent_rdata_fifo|always4~0_combout ),
	.mem_0_0(\data_i_s1_agent_rdata_fifo|mem[0][0]~q ),
	.av_readdata_pre_1(\data_i_s1_translator|av_readdata_pre[1]~q ),
	.mem_1_0(\data_i_s1_agent_rdata_fifo|mem[0][1]~q ),
	.av_readdata_pre_2(\data_i_s1_translator|av_readdata_pre[2]~q ),
	.mem_2_0(\data_i_s1_agent_rdata_fifo|mem[0][2]~q ),
	.av_readdata_pre_3(\data_i_s1_translator|av_readdata_pre[3]~q ),
	.mem_3_0(\data_i_s1_agent_rdata_fifo|mem[0][3]~q ),
	.av_readdata_pre_4(\data_i_s1_translator|av_readdata_pre[4]~q ),
	.mem_4_0(\data_i_s1_agent_rdata_fifo|mem[0][4]~q ),
	.av_readdata_pre_5(\data_i_s1_translator|av_readdata_pre[5]~q ),
	.mem_5_0(\data_i_s1_agent_rdata_fifo|mem[0][5]~q ),
	.av_readdata_pre_6(\data_i_s1_translator|av_readdata_pre[6]~q ),
	.mem_6_0(\data_i_s1_agent_rdata_fifo|mem[0][6]~q ),
	.av_readdata_pre_7(\data_i_s1_translator|av_readdata_pre[7]~q ),
	.mem_7_0(\data_i_s1_agent_rdata_fifo|mem[0][7]~q ),
	.av_readdata_pre_8(\data_i_s1_translator|av_readdata_pre[8]~q ),
	.mem_8_0(\data_i_s1_agent_rdata_fifo|mem[0][8]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.WideOr0(\rsp_demux_005|WideOr0~0_combout ),
	.clk(clk_clk));

spw_babasu_altera_avalon_sc_fifo_5 data_i_s1_agent_rsp_fifo(
	.out_valid_reg(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\data_i_s1_agent_rsp_fifo|mem_used[1]~q ),
	.WideOr0(\data_i_s1_agent|WideOr0~0_combout ),
	.in_data_reg_68(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ),
	.stateST_UNCOMP_WR_SUBBURST(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.mem_129_0(\data_i_s1_agent_rsp_fifo|mem[0][129]~q ),
	.mem_used_0(\data_i_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_68_0(\data_i_s1_agent_rsp_fifo|mem[0][68]~q ),
	.mem_66_0(\data_i_s1_agent_rsp_fifo|mem[0][66]~q ),
	.comb(\data_i_s1_agent|comb~0_combout ),
	.mem_130_0(\data_i_s1_agent_rsp_fifo|mem[0][130]~q ),
	.mem_78_0(\data_i_s1_agent_rsp_fifo|mem[0][78]~q ),
	.mem_77_0(\data_i_s1_agent_rsp_fifo|mem[0][77]~q ),
	.mem_76_0(\data_i_s1_agent_rsp_fifo|mem[0][76]~q ),
	.mem_75_0(\data_i_s1_agent_rsp_fifo|mem[0][75]~q ),
	.mem_74_0(\data_i_s1_agent_rsp_fifo|mem[0][74]~q ),
	.mem_105_0(\data_i_s1_agent_rsp_fifo|mem[0][105]~q ),
	.mem_106_0(\data_i_s1_agent_rsp_fifo|mem[0][106]~q ),
	.mem_107_0(\data_i_s1_agent_rsp_fifo|mem[0][107]~q ),
	.mem_108_0(\data_i_s1_agent_rsp_fifo|mem[0][108]~q ),
	.mem_109_0(\data_i_s1_agent_rsp_fifo|mem[0][109]~q ),
	.mem_110_0(\data_i_s1_agent_rsp_fifo|mem[0][110]~q ),
	.mem_111_0(\data_i_s1_agent_rsp_fifo|mem[0][111]~q ),
	.mem_112_0(\data_i_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_113_0(\data_i_s1_agent_rsp_fifo|mem[0][113]~q ),
	.mem_114_0(\data_i_s1_agent_rsp_fifo|mem[0][114]~q ),
	.mem_115_0(\data_i_s1_agent_rsp_fifo|mem[0][115]~q ),
	.mem_116_0(\data_i_s1_agent_rsp_fifo|mem[0][116]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.nxt_out_eop(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.last_packet_beat(\data_i_s1_agent|uncompressor|last_packet_beat~2_combout ),
	.WideOr01(\rsp_demux_005|WideOr0~0_combout ),
	.read(\data_i_s1_agent_rsp_fifo|read~0_combout ),
	.cp_ready(\data_i_s1_agent|cp_ready~4_combout ),
	.in_data_reg_69(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.rf_source_valid(\data_i_s1_agent|rf_source_valid~0_combout ),
	.out_byte_cnt_reg_2(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_3(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_4(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_5(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_6(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.sink_ready(\data_i_s1_agent|uncompressor|sink_ready~0_combout ),
	.in_data_reg_105(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ),
	.in_data_reg_106(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ),
	.in_data_reg_107(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ),
	.in_data_reg_108(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ),
	.in_data_reg_109(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ),
	.in_data_reg_110(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ),
	.in_data_reg_111(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ),
	.in_data_reg_112(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ),
	.in_data_reg_113(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ),
	.in_data_reg_114(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ),
	.in_data_reg_115(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ),
	.in_data_reg_116(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ),
	.clk(clk_clk));

spw_babasu_altera_avalon_sc_fifo_17 rx_empty_s1_agent_rsp_fifo(
	.h2f_RREADY_0(h2f_RREADY_0),
	.waitrequest_reset_override(\autostart_s1_translator|waitrequest_reset_override~q ),
	.mem_used_1(\rx_empty_s1_agent_rsp_fifo|mem_used[1]~q ),
	.in_data_reg_69(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.wait_latency_counter_1(\rx_empty_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\rx_empty_s1_translator|wait_latency_counter[0]~q ),
	.nxt_out_eop(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.out_valid_reg(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.stateST_UNCOMP_WR_SUBBURST(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.mem_130_0(\rx_empty_s1_agent_rsp_fifo|mem[0][130]~q ),
	.empty(\rx_empty_s1_agent_rdata_fifo|empty~combout ),
	.mem_66_0(\rx_empty_s1_agent_rsp_fifo|mem[0][66]~q ),
	.mem_used_0(\rx_empty_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_78_0(\rx_empty_s1_agent_rsp_fifo|mem[0][78]~q ),
	.mem_77_0(\rx_empty_s1_agent_rsp_fifo|mem[0][77]~q ),
	.mem_76_0(\rx_empty_s1_agent_rsp_fifo|mem[0][76]~q ),
	.mem_75_0(\rx_empty_s1_agent_rsp_fifo|mem[0][75]~q ),
	.mem_74_0(\rx_empty_s1_agent_rsp_fifo|mem[0][74]~q ),
	.mem_105_0(\rx_empty_s1_agent_rsp_fifo|mem[0][105]~q ),
	.mem_106_0(\rx_empty_s1_agent_rsp_fifo|mem[0][106]~q ),
	.mem_107_0(\rx_empty_s1_agent_rsp_fifo|mem[0][107]~q ),
	.mem_108_0(\rx_empty_s1_agent_rsp_fifo|mem[0][108]~q ),
	.mem_109_0(\rx_empty_s1_agent_rsp_fifo|mem[0][109]~q ),
	.mem_110_0(\rx_empty_s1_agent_rsp_fifo|mem[0][110]~q ),
	.mem_111_0(\rx_empty_s1_agent_rsp_fifo|mem[0][111]~q ),
	.mem_112_0(\rx_empty_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_113_0(\rx_empty_s1_agent_rsp_fifo|mem[0][113]~q ),
	.mem_114_0(\rx_empty_s1_agent_rsp_fifo|mem[0][114]~q ),
	.mem_115_0(\rx_empty_s1_agent_rsp_fifo|mem[0][115]~q ),
	.mem_116_0(\rx_empty_s1_agent_rsp_fifo|mem[0][116]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.last_packet_beat(\rx_empty_s1_agent|uncompressor|last_packet_beat~2_combout ),
	.write(\rx_empty_s1_agent_rsp_fifo|write~0_combout ),
	.write1(\rx_empty_s1_agent_rsp_fifo|write~1_combout ),
	.out_byte_cnt_reg_2(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_5(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_4(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_3(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_6(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.in_data_reg_105(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ),
	.in_data_reg_106(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ),
	.in_data_reg_107(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ),
	.in_data_reg_108(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ),
	.in_data_reg_109(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ),
	.in_data_reg_110(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ),
	.in_data_reg_111(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ),
	.in_data_reg_112(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ),
	.in_data_reg_113(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ),
	.in_data_reg_114(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ),
	.in_data_reg_115(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ),
	.in_data_reg_116(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ),
	.clk(clk_clk));

spw_babasu_altera_merlin_slave_agent_8 rx_empty_s1_agent(
	.h2f_RREADY_0(h2f_RREADY_0),
	.waitrequest_reset_override(\autostart_s1_translator|waitrequest_reset_override~q ),
	.stateST_COMP_TRANS(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.mem_used_1(\rx_empty_s1_agent_rsp_fifo|mem_used[1]~q ),
	.in_data_reg_69(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.in_narrow_reg(\rx_empty_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.wait_latency_counter_1(\rx_empty_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\rx_empty_s1_translator|wait_latency_counter[0]~q ),
	.cp_ready(\rx_empty_s1_agent|cp_ready~0_combout ),
	.cp_ready1(\rx_empty_s1_agent|cp_ready~1_combout ),
	.empty(\rx_empty_s1_agent_rdata_fifo|empty~combout ),
	.mem_66_0(\rx_empty_s1_agent_rsp_fifo|mem[0][66]~q ),
	.mem_used_0(\rx_empty_s1_agent_rsp_fifo|mem_used[0]~q ),
	.last_packet_beat(\rx_empty_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.mem_78_0(\rx_empty_s1_agent_rsp_fifo|mem[0][78]~q ),
	.mem_77_0(\rx_empty_s1_agent_rsp_fifo|mem[0][77]~q ),
	.mem_76_0(\rx_empty_s1_agent_rsp_fifo|mem[0][76]~q ),
	.mem_75_0(\rx_empty_s1_agent_rsp_fifo|mem[0][75]~q ),
	.mem_74_0(\rx_empty_s1_agent_rsp_fifo|mem[0][74]~q ),
	.last_packet_beat1(\rx_empty_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.last_packet_beat2(\rx_empty_s1_agent|uncompressor|last_packet_beat~2_combout ),
	.cp_ready2(\rx_empty_s1_agent|cp_ready~2_combout ),
	.clk_clk(clk_clk));

spw_babasu_altera_avalon_sc_fifo_14 rd_data_s1_agent_rdata_fifo(
	.read_latency_shift_reg_0(\rd_data_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\rd_data_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_129_0(\rd_data_s1_agent_rsp_fifo|mem[0][129]~q ),
	.mem_used_01(\rd_data_s1_agent_rsp_fifo|mem_used[0]~q ),
	.av_readdata_pre_0(\rd_data_s1_translator|av_readdata_pre[0]~q ),
	.mem_0_0(\rd_data_s1_agent_rdata_fifo|mem[0][0]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.WideOr0(\rsp_demux_009|WideOr0~0_combout ),
	.clk(clk_clk));

spw_babasu_altera_avalon_sc_fifo_15 rd_data_s1_agent_rsp_fifo(
	.out_valid_reg(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\rd_data_s1_agent_rsp_fifo|mem_used[1]~q ),
	.WideOr0(\rd_data_s1_agent|WideOr0~0_combout ),
	.in_data_reg_68(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ),
	.stateST_UNCOMP_WR_SUBBURST(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.mem_129_0(\rd_data_s1_agent_rsp_fifo|mem[0][129]~q ),
	.mem_used_0(\rd_data_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_68_0(\rd_data_s1_agent_rsp_fifo|mem[0][68]~q ),
	.mem_66_0(\rd_data_s1_agent_rsp_fifo|mem[0][66]~q ),
	.comb(\rd_data_s1_agent|comb~0_combout ),
	.mem_130_0(\rd_data_s1_agent_rsp_fifo|mem[0][130]~q ),
	.mem_78_0(\rd_data_s1_agent_rsp_fifo|mem[0][78]~q ),
	.mem_77_0(\rd_data_s1_agent_rsp_fifo|mem[0][77]~q ),
	.mem_76_0(\rd_data_s1_agent_rsp_fifo|mem[0][76]~q ),
	.mem_75_0(\rd_data_s1_agent_rsp_fifo|mem[0][75]~q ),
	.mem_74_0(\rd_data_s1_agent_rsp_fifo|mem[0][74]~q ),
	.mem_105_0(\rd_data_s1_agent_rsp_fifo|mem[0][105]~q ),
	.mem_106_0(\rd_data_s1_agent_rsp_fifo|mem[0][106]~q ),
	.mem_107_0(\rd_data_s1_agent_rsp_fifo|mem[0][107]~q ),
	.mem_108_0(\rd_data_s1_agent_rsp_fifo|mem[0][108]~q ),
	.mem_109_0(\rd_data_s1_agent_rsp_fifo|mem[0][109]~q ),
	.mem_110_0(\rd_data_s1_agent_rsp_fifo|mem[0][110]~q ),
	.mem_111_0(\rd_data_s1_agent_rsp_fifo|mem[0][111]~q ),
	.mem_112_0(\rd_data_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_113_0(\rd_data_s1_agent_rsp_fifo|mem[0][113]~q ),
	.mem_114_0(\rd_data_s1_agent_rsp_fifo|mem[0][114]~q ),
	.mem_115_0(\rd_data_s1_agent_rsp_fifo|mem[0][115]~q ),
	.mem_116_0(\rd_data_s1_agent_rsp_fifo|mem[0][116]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.nxt_out_eop(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.last_packet_beat(\rd_data_s1_agent|uncompressor|last_packet_beat~2_combout ),
	.WideOr01(\rsp_demux_009|WideOr0~0_combout ),
	.read(\rd_data_s1_agent_rsp_fifo|read~0_combout ),
	.cp_ready(\rd_data_s1_agent|cp_ready~4_combout ),
	.in_data_reg_69(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.rf_source_valid(\rd_data_s1_agent|rf_source_valid~0_combout ),
	.out_byte_cnt_reg_2(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_4(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_3(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_5(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_6(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.sink_ready(\rd_data_s1_agent|uncompressor|sink_ready~0_combout ),
	.in_data_reg_105(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ),
	.in_data_reg_106(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ),
	.in_data_reg_107(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ),
	.in_data_reg_108(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ),
	.in_data_reg_109(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ),
	.in_data_reg_110(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ),
	.in_data_reg_111(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ),
	.in_data_reg_112(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ),
	.in_data_reg_113(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ),
	.in_data_reg_114(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ),
	.in_data_reg_115(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ),
	.in_data_reg_116(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ),
	.clk(clk_clk));

spw_babasu_altera_merlin_slave_agent_7 rd_data_s1_agent(
	.waitrequest_reset_override(\autostart_s1_translator|waitrequest_reset_override~q ),
	.stateST_COMP_TRANS(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.out_valid_reg(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\rd_data_s1_agent_rsp_fifo|mem_used[1]~q ),
	.in_narrow_reg(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.in_byteen_reg_3(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ),
	.in_byteen_reg_2(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ),
	.in_byteen_reg_1(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ),
	.in_byteen_reg_0(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ),
	.WideOr0(\rd_data_s1_agent|WideOr0~0_combout ),
	.wait_latency_counter_1(wait_latency_counter_16),
	.wait_latency_counter_0(wait_latency_counter_06),
	.in_data_reg_68(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ),
	.cp_ready(\rd_data_s1_agent|cp_ready~0_combout ),
	.read_latency_shift_reg_0(\rd_data_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\rd_data_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_129_0(\rd_data_s1_agent_rsp_fifo|mem[0][129]~q ),
	.mem_used_01(\rd_data_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_66_0(\rd_data_s1_agent_rsp_fifo|mem[0][66]~q ),
	.comb(\rd_data_s1_agent|comb~0_combout ),
	.last_packet_beat(\rd_data_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.mem_78_0(\rd_data_s1_agent_rsp_fifo|mem[0][78]~q ),
	.mem_77_0(\rd_data_s1_agent_rsp_fifo|mem[0][77]~q ),
	.mem_76_0(\rd_data_s1_agent_rsp_fifo|mem[0][76]~q ),
	.mem_75_0(\rd_data_s1_agent_rsp_fifo|mem[0][75]~q ),
	.mem_74_0(\rd_data_s1_agent_rsp_fifo|mem[0][74]~q ),
	.last_packet_beat1(\rd_data_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.m0_write1(m0_write4),
	.nxt_out_eop(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.cp_ready1(\rd_data_s1_agent|cp_ready~3_combout ),
	.last_packet_beat2(\rd_data_s1_agent|uncompressor|last_packet_beat~2_combout ),
	.WideOr01(\rsp_demux_009|WideOr0~0_combout ),
	.read(\rd_data_s1_agent_rsp_fifo|read~0_combout ),
	.cp_ready2(\rd_data_s1_agent|cp_ready~4_combout ),
	.in_data_reg_69(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.rf_source_valid(\rd_data_s1_agent|rf_source_valid~0_combout ),
	.rf_sink_ready(\rd_data_s1_agent|uncompressor|sink_ready~0_combout ),
	.clk_clk(clk_clk));

spw_babasu_altera_avalon_sc_fifo_6 data_o_s1_agent_rdata_fifo(
	.h2f_RREADY_0(h2f_RREADY_0),
	.read_latency_shift_reg_0(\data_o_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\data_o_s1_agent_rdata_fifo|mem_used[0]~q ),
	.empty1(\data_o_s1_agent_rdata_fifo|empty~combout ),
	.av_readdata_pre_0(\data_o_s1_translator|av_readdata_pre[0]~q ),
	.mem_0_0(\data_o_s1_agent_rdata_fifo|mem[0][0]~q ),
	.mem_1_0(\data_o_s1_agent_rdata_fifo|mem[0][1]~q ),
	.av_readdata_pre_1(\data_o_s1_translator|av_readdata_pre[1]~q ),
	.mem_2_0(\data_o_s1_agent_rdata_fifo|mem[0][2]~q ),
	.av_readdata_pre_2(\data_o_s1_translator|av_readdata_pre[2]~q ),
	.mem_3_0(\data_o_s1_agent_rdata_fifo|mem[0][3]~q ),
	.av_readdata_pre_3(\data_o_s1_translator|av_readdata_pre[3]~q ),
	.mem_4_0(\data_o_s1_agent_rdata_fifo|mem[0][4]~q ),
	.av_readdata_pre_4(\data_o_s1_translator|av_readdata_pre[4]~q ),
	.mem_5_0(\data_o_s1_agent_rdata_fifo|mem[0][5]~q ),
	.av_readdata_pre_5(\data_o_s1_translator|av_readdata_pre[5]~q ),
	.mem_6_0(\data_o_s1_agent_rdata_fifo|mem[0][6]~q ),
	.av_readdata_pre_6(\data_o_s1_translator|av_readdata_pre[6]~q ),
	.mem_7_0(\data_o_s1_agent_rdata_fifo|mem[0][7]~q ),
	.av_readdata_pre_7(\data_o_s1_translator|av_readdata_pre[7]~q ),
	.mem_8_0(\data_o_s1_agent_rdata_fifo|mem[0][8]~q ),
	.av_readdata_pre_8(\data_o_s1_translator|av_readdata_pre[8]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.clk(clk_clk));

spw_babasu_altera_avalon_sc_fifo_7 data_o_s1_agent_rsp_fifo(
	.h2f_RREADY_0(h2f_RREADY_0),
	.mem_used_1(\data_o_s1_agent_rsp_fifo|mem_used[1]~q ),
	.waitrequest_reset_override(\autostart_s1_translator|waitrequest_reset_override~q ),
	.in_data_reg_69(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.wait_latency_counter_1(\data_o_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\data_o_s1_translator|wait_latency_counter[0]~q ),
	.nxt_out_eop(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.out_valid_reg(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.stateST_UNCOMP_WR_SUBBURST(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.mem_130_0(\data_o_s1_agent_rsp_fifo|mem[0][130]~q ),
	.empty(\data_o_s1_agent_rdata_fifo|empty~combout ),
	.mem_66_0(\data_o_s1_agent_rsp_fifo|mem[0][66]~q ),
	.mem_used_0(\data_o_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_78_0(\data_o_s1_agent_rsp_fifo|mem[0][78]~q ),
	.mem_77_0(\data_o_s1_agent_rsp_fifo|mem[0][77]~q ),
	.mem_76_0(\data_o_s1_agent_rsp_fifo|mem[0][76]~q ),
	.mem_75_0(\data_o_s1_agent_rsp_fifo|mem[0][75]~q ),
	.mem_74_0(\data_o_s1_agent_rsp_fifo|mem[0][74]~q ),
	.mem_105_0(\data_o_s1_agent_rsp_fifo|mem[0][105]~q ),
	.mem_106_0(\data_o_s1_agent_rsp_fifo|mem[0][106]~q ),
	.mem_107_0(\data_o_s1_agent_rsp_fifo|mem[0][107]~q ),
	.mem_108_0(\data_o_s1_agent_rsp_fifo|mem[0][108]~q ),
	.mem_109_0(\data_o_s1_agent_rsp_fifo|mem[0][109]~q ),
	.mem_110_0(\data_o_s1_agent_rsp_fifo|mem[0][110]~q ),
	.mem_111_0(\data_o_s1_agent_rsp_fifo|mem[0][111]~q ),
	.mem_112_0(\data_o_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_113_0(\data_o_s1_agent_rsp_fifo|mem[0][113]~q ),
	.mem_114_0(\data_o_s1_agent_rsp_fifo|mem[0][114]~q ),
	.mem_115_0(\data_o_s1_agent_rsp_fifo|mem[0][115]~q ),
	.mem_116_0(\data_o_s1_agent_rsp_fifo|mem[0][116]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.last_packet_beat(\data_o_s1_agent|uncompressor|last_packet_beat~2_combout ),
	.write(\data_o_s1_agent_rsp_fifo|write~0_combout ),
	.write1(\data_o_s1_agent_rsp_fifo|write~1_combout ),
	.out_byte_cnt_reg_2(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_6(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.out_uncomp_byte_cnt_reg_5(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_4(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_3(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.in_data_reg_105(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ),
	.in_data_reg_106(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ),
	.in_data_reg_107(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ),
	.in_data_reg_108(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ),
	.in_data_reg_109(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ),
	.in_data_reg_110(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ),
	.in_data_reg_111(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ),
	.in_data_reg_112(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ),
	.in_data_reg_113(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ),
	.in_data_reg_114(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ),
	.in_data_reg_115(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ),
	.in_data_reg_116(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ),
	.clk(clk_clk));

spw_babasu_altera_merlin_slave_agent_3 data_o_s1_agent(
	.h2f_RREADY_0(h2f_RREADY_0),
	.stateST_COMP_TRANS(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.mem_used_1(\data_o_s1_agent_rsp_fifo|mem_used[1]~q ),
	.waitrequest_reset_override(\autostart_s1_translator|waitrequest_reset_override~q ),
	.in_data_reg_69(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.in_narrow_reg(\data_o_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.wait_latency_counter_1(\data_o_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\data_o_s1_translator|wait_latency_counter[0]~q ),
	.cp_ready(\data_o_s1_agent|cp_ready~0_combout ),
	.cp_ready1(\data_o_s1_agent|cp_ready~1_combout ),
	.empty(\data_o_s1_agent_rdata_fifo|empty~combout ),
	.mem_66_0(\data_o_s1_agent_rsp_fifo|mem[0][66]~q ),
	.mem_used_0(\data_o_s1_agent_rsp_fifo|mem_used[0]~q ),
	.last_packet_beat(\data_o_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.mem_78_0(\data_o_s1_agent_rsp_fifo|mem[0][78]~q ),
	.mem_77_0(\data_o_s1_agent_rsp_fifo|mem[0][77]~q ),
	.mem_76_0(\data_o_s1_agent_rsp_fifo|mem[0][76]~q ),
	.mem_75_0(\data_o_s1_agent_rsp_fifo|mem[0][75]~q ),
	.mem_74_0(\data_o_s1_agent_rsp_fifo|mem[0][74]~q ),
	.last_packet_beat1(\data_o_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.last_packet_beat2(\data_o_s1_agent|uncompressor|last_packet_beat~2_combout ),
	.cp_ready2(\data_o_s1_agent|cp_ready~2_combout ),
	.clk_clk(clk_clk));

spw_babasu_altera_avalon_sc_fifo_30 tx_full_s1_agent_rdata_fifo(
	.h2f_RREADY_0(h2f_RREADY_0),
	.read_latency_shift_reg_0(\tx_full_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\tx_full_s1_agent_rdata_fifo|mem_used[0]~q ),
	.empty1(\tx_full_s1_agent_rdata_fifo|empty~combout ),
	.mem_0_0(\tx_full_s1_agent_rdata_fifo|mem[0][0]~q ),
	.av_readdata_pre_0(\tx_full_s1_translator|av_readdata_pre[0]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.clk(clk_clk));

spw_babasu_altera_avalon_sc_fifo_31 tx_full_s1_agent_rsp_fifo(
	.h2f_RREADY_0(h2f_RREADY_0),
	.waitrequest_reset_override(\autostart_s1_translator|waitrequest_reset_override~q ),
	.in_data_reg_69(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.mem_used_1(\tx_full_s1_agent_rsp_fifo|mem_used[1]~q ),
	.wait_latency_counter_1(\tx_full_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\tx_full_s1_translator|wait_latency_counter[0]~q ),
	.out_valid_reg(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.stateST_UNCOMP_WR_SUBBURST(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.empty(\tx_full_s1_agent_rdata_fifo|empty~combout ),
	.mem_66_0(\tx_full_s1_agent_rsp_fifo|mem[0][66]~q ),
	.mem_used_0(\tx_full_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_78_0(\tx_full_s1_agent_rsp_fifo|mem[0][78]~q ),
	.mem_77_0(\tx_full_s1_agent_rsp_fifo|mem[0][77]~q ),
	.mem_76_0(\tx_full_s1_agent_rsp_fifo|mem[0][76]~q ),
	.mem_75_0(\tx_full_s1_agent_rsp_fifo|mem[0][75]~q ),
	.mem_74_0(\tx_full_s1_agent_rsp_fifo|mem[0][74]~q ),
	.last_packet_beat(\tx_full_s1_agent|uncompressor|last_packet_beat~3_combout ),
	.mem_130_0(\tx_full_s1_agent_rsp_fifo|mem[0][130]~q ),
	.mem_105_0(\tx_full_s1_agent_rsp_fifo|mem[0][105]~q ),
	.mem_106_0(\tx_full_s1_agent_rsp_fifo|mem[0][106]~q ),
	.mem_107_0(\tx_full_s1_agent_rsp_fifo|mem[0][107]~q ),
	.mem_108_0(\tx_full_s1_agent_rsp_fifo|mem[0][108]~q ),
	.mem_109_0(\tx_full_s1_agent_rsp_fifo|mem[0][109]~q ),
	.mem_110_0(\tx_full_s1_agent_rsp_fifo|mem[0][110]~q ),
	.mem_111_0(\tx_full_s1_agent_rsp_fifo|mem[0][111]~q ),
	.mem_112_0(\tx_full_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_113_0(\tx_full_s1_agent_rsp_fifo|mem[0][113]~q ),
	.mem_114_0(\tx_full_s1_agent_rsp_fifo|mem[0][114]~q ),
	.mem_115_0(\tx_full_s1_agent_rsp_fifo|mem[0][115]~q ),
	.mem_116_0(\tx_full_s1_agent_rsp_fifo|mem[0][116]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.nxt_out_eop(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.out_byte_cnt_reg_2(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.write(\tx_full_s1_agent_rsp_fifo|write~0_combout ),
	.write1(\tx_full_s1_agent_rsp_fifo|write~1_combout ),
	.out_uncomp_byte_cnt_reg_3(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_6(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.out_uncomp_byte_cnt_reg_5(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_4(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.in_data_reg_105(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ),
	.in_data_reg_106(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ),
	.in_data_reg_107(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ),
	.in_data_reg_108(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ),
	.in_data_reg_109(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ),
	.in_data_reg_110(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ),
	.in_data_reg_111(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ),
	.in_data_reg_112(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ),
	.in_data_reg_113(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ),
	.in_data_reg_114(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ),
	.in_data_reg_115(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ),
	.in_data_reg_116(\tx_full_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ),
	.clk(clk_clk));

spw_babasu_altera_avalon_sc_fifo_11 link_disable_s1_agent_rsp_fifo(
	.out_valid_reg(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\link_disable_s1_agent_rsp_fifo|mem_used[1]~q ),
	.WideOr0(\link_disable_s1_agent|WideOr0~0_combout ),
	.in_data_reg_68(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ),
	.stateST_UNCOMP_WR_SUBBURST(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.mem_129_0(\link_disable_s1_agent_rsp_fifo|mem[0][129]~q ),
	.mem_used_0(\link_disable_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_68_0(\link_disable_s1_agent_rsp_fifo|mem[0][68]~q ),
	.mem_66_0(\link_disable_s1_agent_rsp_fifo|mem[0][66]~q ),
	.comb(\link_disable_s1_agent|comb~0_combout ),
	.mem_130_0(\link_disable_s1_agent_rsp_fifo|mem[0][130]~q ),
	.mem_78_0(\link_disable_s1_agent_rsp_fifo|mem[0][78]~q ),
	.mem_77_0(\link_disable_s1_agent_rsp_fifo|mem[0][77]~q ),
	.mem_76_0(\link_disable_s1_agent_rsp_fifo|mem[0][76]~q ),
	.mem_75_0(\link_disable_s1_agent_rsp_fifo|mem[0][75]~q ),
	.mem_74_0(\link_disable_s1_agent_rsp_fifo|mem[0][74]~q ),
	.mem_105_0(\link_disable_s1_agent_rsp_fifo|mem[0][105]~q ),
	.mem_106_0(\link_disable_s1_agent_rsp_fifo|mem[0][106]~q ),
	.mem_107_0(\link_disable_s1_agent_rsp_fifo|mem[0][107]~q ),
	.mem_108_0(\link_disable_s1_agent_rsp_fifo|mem[0][108]~q ),
	.mem_109_0(\link_disable_s1_agent_rsp_fifo|mem[0][109]~q ),
	.mem_110_0(\link_disable_s1_agent_rsp_fifo|mem[0][110]~q ),
	.mem_111_0(\link_disable_s1_agent_rsp_fifo|mem[0][111]~q ),
	.mem_112_0(\link_disable_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_113_0(\link_disable_s1_agent_rsp_fifo|mem[0][113]~q ),
	.mem_114_0(\link_disable_s1_agent_rsp_fifo|mem[0][114]~q ),
	.mem_115_0(\link_disable_s1_agent_rsp_fifo|mem[0][115]~q ),
	.mem_116_0(\link_disable_s1_agent_rsp_fifo|mem[0][116]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.nxt_out_eop(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.last_packet_beat(\link_disable_s1_agent|uncompressor|last_packet_beat~2_combout ),
	.WideOr01(\rsp_demux_001|WideOr0~0_combout ),
	.read(\link_disable_s1_agent_rsp_fifo|read~0_combout ),
	.cp_ready(\link_disable_s1_agent|cp_ready~4_combout ),
	.in_data_reg_69(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.rf_source_valid(\link_disable_s1_agent|rf_source_valid~0_combout ),
	.out_byte_cnt_reg_2(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_3(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_4(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_5(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_6(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.sink_ready(\link_disable_s1_agent|uncompressor|sink_ready~0_combout ),
	.in_data_reg_105(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ),
	.in_data_reg_106(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ),
	.in_data_reg_107(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ),
	.in_data_reg_108(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ),
	.in_data_reg_109(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ),
	.in_data_reg_110(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ),
	.in_data_reg_111(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ),
	.in_data_reg_112(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ),
	.in_data_reg_113(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ),
	.in_data_reg_114(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ),
	.in_data_reg_115(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ),
	.in_data_reg_116(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ),
	.clk(clk_clk));

spw_babasu_altera_merlin_slave_agent_5 link_disable_s1_agent(
	.waitrequest_reset_override(\autostart_s1_translator|waitrequest_reset_override~q ),
	.stateST_COMP_TRANS(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.out_valid_reg(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\link_disable_s1_agent_rsp_fifo|mem_used[1]~q ),
	.in_narrow_reg(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.in_byteen_reg_3(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ),
	.in_byteen_reg_2(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ),
	.in_byteen_reg_1(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ),
	.in_byteen_reg_0(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ),
	.WideOr0(\link_disable_s1_agent|WideOr0~0_combout ),
	.wait_latency_counter_1(wait_latency_counter_1),
	.wait_latency_counter_0(wait_latency_counter_0),
	.in_data_reg_68(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ),
	.cp_ready(\link_disable_s1_agent|cp_ready~0_combout ),
	.read_latency_shift_reg_0(\link_disable_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\link_disable_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_129_0(\link_disable_s1_agent_rsp_fifo|mem[0][129]~q ),
	.mem_used_01(\link_disable_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_66_0(\link_disable_s1_agent_rsp_fifo|mem[0][66]~q ),
	.comb(\link_disable_s1_agent|comb~0_combout ),
	.last_packet_beat(\link_disable_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.mem_78_0(\link_disable_s1_agent_rsp_fifo|mem[0][78]~q ),
	.mem_77_0(\link_disable_s1_agent_rsp_fifo|mem[0][77]~q ),
	.mem_76_0(\link_disable_s1_agent_rsp_fifo|mem[0][76]~q ),
	.mem_75_0(\link_disable_s1_agent_rsp_fifo|mem[0][75]~q ),
	.mem_74_0(\link_disable_s1_agent_rsp_fifo|mem[0][74]~q ),
	.last_packet_beat1(\link_disable_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.m0_write1(m0_write2),
	.nxt_out_eop(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.cp_ready1(\link_disable_s1_agent|cp_ready~3_combout ),
	.last_packet_beat2(\link_disable_s1_agent|uncompressor|last_packet_beat~2_combout ),
	.WideOr01(\rsp_demux_001|WideOr0~0_combout ),
	.read(\link_disable_s1_agent_rsp_fifo|read~0_combout ),
	.cp_ready2(\link_disable_s1_agent|cp_ready~4_combout ),
	.in_data_reg_69(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.rf_source_valid(\link_disable_s1_agent|rf_source_valid~0_combout ),
	.rf_sink_ready(\link_disable_s1_agent|uncompressor|sink_ready~0_combout ),
	.clk_clk(clk_clk));

spw_babasu_altera_avalon_sc_fifo_12 link_start_s1_agent_rdata_fifo(
	.read_latency_shift_reg_0(\link_start_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\link_start_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_129_0(\link_start_s1_agent_rsp_fifo|mem[0][129]~q ),
	.mem_used_01(\link_start_s1_agent_rsp_fifo|mem_used[0]~q ),
	.av_readdata_pre_0(\link_start_s1_translator|av_readdata_pre[0]~q ),
	.mem_0_0(\link_start_s1_agent_rdata_fifo|mem[0][0]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.WideOr0(\rsp_demux|WideOr0~0_combout ),
	.clk(clk_clk));

spw_babasu_altera_avalon_sc_fifo_13 link_start_s1_agent_rsp_fifo(
	.out_valid_reg(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\link_start_s1_agent_rsp_fifo|mem_used[1]~q ),
	.WideOr0(\link_start_s1_agent|WideOr0~0_combout ),
	.in_data_reg_68(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ),
	.stateST_UNCOMP_WR_SUBBURST(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.mem_129_0(\link_start_s1_agent_rsp_fifo|mem[0][129]~q ),
	.mem_used_0(\link_start_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_68_0(\link_start_s1_agent_rsp_fifo|mem[0][68]~q ),
	.mem_66_0(\link_start_s1_agent_rsp_fifo|mem[0][66]~q ),
	.comb(\link_start_s1_agent|comb~0_combout ),
	.mem_130_0(\link_start_s1_agent_rsp_fifo|mem[0][130]~q ),
	.mem_78_0(\link_start_s1_agent_rsp_fifo|mem[0][78]~q ),
	.mem_77_0(\link_start_s1_agent_rsp_fifo|mem[0][77]~q ),
	.mem_76_0(\link_start_s1_agent_rsp_fifo|mem[0][76]~q ),
	.mem_75_0(\link_start_s1_agent_rsp_fifo|mem[0][75]~q ),
	.mem_74_0(\link_start_s1_agent_rsp_fifo|mem[0][74]~q ),
	.mem_105_0(\link_start_s1_agent_rsp_fifo|mem[0][105]~q ),
	.mem_106_0(\link_start_s1_agent_rsp_fifo|mem[0][106]~q ),
	.mem_107_0(\link_start_s1_agent_rsp_fifo|mem[0][107]~q ),
	.mem_108_0(\link_start_s1_agent_rsp_fifo|mem[0][108]~q ),
	.mem_109_0(\link_start_s1_agent_rsp_fifo|mem[0][109]~q ),
	.mem_110_0(\link_start_s1_agent_rsp_fifo|mem[0][110]~q ),
	.mem_111_0(\link_start_s1_agent_rsp_fifo|mem[0][111]~q ),
	.mem_112_0(\link_start_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_113_0(\link_start_s1_agent_rsp_fifo|mem[0][113]~q ),
	.mem_114_0(\link_start_s1_agent_rsp_fifo|mem[0][114]~q ),
	.mem_115_0(\link_start_s1_agent_rsp_fifo|mem[0][115]~q ),
	.mem_116_0(\link_start_s1_agent_rsp_fifo|mem[0][116]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.nxt_out_eop(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.last_packet_beat(\link_start_s1_agent|uncompressor|last_packet_beat~2_combout ),
	.WideOr01(\rsp_demux|WideOr0~0_combout ),
	.read(\link_start_s1_agent_rsp_fifo|read~0_combout ),
	.cp_ready(\link_start_s1_agent|cp_ready~3_combout ),
	.in_data_reg_69(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.rf_source_valid(\link_start_s1_agent|rf_source_valid~0_combout ),
	.out_byte_cnt_reg_2(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_3(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_4(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_5(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_6(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.sink_ready(\link_start_s1_agent|uncompressor|sink_ready~0_combout ),
	.in_data_reg_105(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ),
	.in_data_reg_106(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ),
	.in_data_reg_107(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ),
	.in_data_reg_108(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ),
	.in_data_reg_109(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ),
	.in_data_reg_110(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ),
	.in_data_reg_111(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ),
	.in_data_reg_112(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ),
	.in_data_reg_113(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[113]~q ),
	.in_data_reg_114(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[114]~q ),
	.in_data_reg_115(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[115]~q ),
	.in_data_reg_116(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[116]~q ),
	.clk(clk_clk));

spw_babasu_altera_merlin_slave_agent_6 link_start_s1_agent(
	.waitrequest_reset_override(\autostart_s1_translator|waitrequest_reset_override~q ),
	.stateST_COMP_TRANS(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.out_valid_reg(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\link_start_s1_agent_rsp_fifo|mem_used[1]~q ),
	.in_narrow_reg(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.in_byteen_reg_3(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ),
	.in_byteen_reg_2(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ),
	.in_byteen_reg_1(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ),
	.in_byteen_reg_0(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ),
	.WideOr0(\link_start_s1_agent|WideOr0~0_combout ),
	.wait_latency_counter_1(wait_latency_counter_17),
	.wait_latency_counter_0(wait_latency_counter_07),
	.in_data_reg_68(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ),
	.cp_ready(\link_start_s1_agent|cp_ready~0_combout ),
	.read_latency_shift_reg_0(\link_start_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\link_start_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_129_0(\link_start_s1_agent_rsp_fifo|mem[0][129]~q ),
	.mem_used_01(\link_start_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_66_0(\link_start_s1_agent_rsp_fifo|mem[0][66]~q ),
	.comb(\link_start_s1_agent|comb~0_combout ),
	.last_packet_beat(\link_start_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.mem_78_0(\link_start_s1_agent_rsp_fifo|mem[0][78]~q ),
	.mem_77_0(\link_start_s1_agent_rsp_fifo|mem[0][77]~q ),
	.mem_76_0(\link_start_s1_agent_rsp_fifo|mem[0][76]~q ),
	.mem_75_0(\link_start_s1_agent_rsp_fifo|mem[0][75]~q ),
	.mem_74_0(\link_start_s1_agent_rsp_fifo|mem[0][74]~q ),
	.last_packet_beat1(\link_start_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.m0_write1(m0_write3),
	.nxt_out_eop(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.cp_ready1(\link_start_s1_agent|cp_ready~2_combout ),
	.last_packet_beat2(\link_start_s1_agent|uncompressor|last_packet_beat~2_combout ),
	.WideOr01(\rsp_demux|WideOr0~0_combout ),
	.read(\link_start_s1_agent_rsp_fifo|read~0_combout ),
	.cp_ready2(\link_start_s1_agent|cp_ready~3_combout ),
	.in_data_reg_69(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.rf_source_valid(\link_start_s1_agent|rf_source_valid~0_combout ),
	.rf_sink_ready(\link_start_s1_agent|uncompressor|sink_ready~0_combout ),
	.clk_clk(clk_clk));

spw_babasu_altera_merlin_axi_master_ni hps_0_h2f_axi_master_agent(
	.h2f_AWVALID_0(h2f_AWVALID_0),
	.h2f_WLAST_0(h2f_WLAST_0),
	.h2f_WVALID_0(h2f_WVALID_0),
	.h2f_ARBURST_0(h2f_ARBURST_0),
	.h2f_ARBURST_1(h2f_ARBURST_1),
	.h2f_ARLEN_0(h2f_ARLEN_0),
	.h2f_ARLEN_1(h2f_ARLEN_1),
	.h2f_ARLEN_2(h2f_ARLEN_2),
	.h2f_ARLEN_3(h2f_ARLEN_3),
	.h2f_ARSIZE_0(h2f_ARSIZE_0),
	.h2f_ARSIZE_1(h2f_ARSIZE_1),
	.h2f_ARSIZE_2(h2f_ARSIZE_2),
	.h2f_AWADDR_0(h2f_AWADDR_0),
	.h2f_AWADDR_1(h2f_AWADDR_1),
	.h2f_AWADDR_2(h2f_AWADDR_2),
	.h2f_AWADDR_3(h2f_AWADDR_3),
	.h2f_AWADDR_4(h2f_AWADDR_4),
	.h2f_AWADDR_5(h2f_AWADDR_5),
	.h2f_AWADDR_6(h2f_AWADDR_6),
	.h2f_AWADDR_7(h2f_AWADDR_7),
	.h2f_AWADDR_8(h2f_AWADDR_8),
	.h2f_AWBURST_0(h2f_AWBURST_0),
	.h2f_AWBURST_1(h2f_AWBURST_1),
	.h2f_AWLEN_0(h2f_AWLEN_0),
	.h2f_AWLEN_1(h2f_AWLEN_1),
	.h2f_AWLEN_2(h2f_AWLEN_2),
	.h2f_AWLEN_3(h2f_AWLEN_3),
	.h2f_AWSIZE_0(h2f_AWSIZE_0),
	.h2f_AWSIZE_1(h2f_AWSIZE_1),
	.h2f_AWSIZE_2(h2f_AWSIZE_2),
	.address_burst_8(\hps_0_h2f_axi_master_agent|align_address_to_size|address_burst[8]~q ),
	.address_burst_7(\hps_0_h2f_axi_master_agent|align_address_to_size|address_burst[7]~q ),
	.address_burst_6(\hps_0_h2f_axi_master_agent|align_address_to_size|address_burst[6]~q ),
	.Add5(\hps_0_h2f_axi_master_agent|Add5~1_sumout ),
	.Add51(\hps_0_h2f_axi_master_agent|Add5~5_sumout ),
	.Add52(\hps_0_h2f_axi_master_agent|Add5~9_sumout ),
	.write_addr_data_both_valid1(\hps_0_h2f_axi_master_agent|write_addr_data_both_valid~combout ),
	.sop_enable1(\hps_0_h2f_axi_master_agent|sop_enable~q ),
	.out_data_8(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[8]~0_combout ),
	.address_burst_5(\hps_0_h2f_axi_master_agent|align_address_to_size|address_burst[5]~q ),
	.out_data_5(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[5]~1_combout ),
	.address_burst_4(\hps_0_h2f_axi_master_agent|align_address_to_size|address_burst[4]~q ),
	.out_data_4(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[4]~2_combout ),
	.out_data_7(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[7]~3_combout ),
	.out_data_6(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[6]~4_combout ),
	.nonposted_cmd_accepted(nonposted_cmd_accepted1),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out1),
	.Decoder1(\hps_0_h2f_axi_master_agent|Decoder1~0_combout ),
	.Add2(\hps_0_h2f_axi_master_agent|Add2~0_combout ),
	.Add21(\hps_0_h2f_axi_master_agent|Add2~1_combout ),
	.Add22(\hps_0_h2f_axi_master_agent|Add2~2_combout ),
	.Add23(\hps_0_h2f_axi_master_agent|Add2~3_combout ),
	.burst_bytecount_5(\hps_0_h2f_axi_master_agent|burst_bytecount[5]~q ),
	.write_cp_data_77(\hps_0_h2f_axi_master_agent|write_cp_data[77]~0_combout ),
	.burst_bytecount_6(\hps_0_h2f_axi_master_agent|burst_bytecount[6]~q ),
	.write_cp_data_78(\hps_0_h2f_axi_master_agent|write_cp_data[78]~1_combout ),
	.burst_bytecount_3(\hps_0_h2f_axi_master_agent|burst_bytecount[3]~q ),
	.write_cp_data_75(\hps_0_h2f_axi_master_agent|write_cp_data[75]~2_combout ),
	.burst_bytecount_2(\hps_0_h2f_axi_master_agent|burst_bytecount[2]~q ),
	.write_cp_data_74(\hps_0_h2f_axi_master_agent|write_cp_data[74]~3_combout ),
	.burst_bytecount_4(\hps_0_h2f_axi_master_agent|burst_bytecount[4]~q ),
	.write_cp_data_76(\hps_0_h2f_axi_master_agent|write_cp_data[76]~4_combout ),
	.Selector3(\hps_0_h2f_axi_master_agent|Selector3~0_combout ),
	.Selector10(\hps_0_h2f_axi_master_agent|Selector10~0_combout ),
	.Selector101(\hps_0_h2f_axi_master_agent|Selector10~1_combout ),
	.base_address_3(\hps_0_h2f_axi_master_agent|align_address_to_size|base_address[3]~0_combout ),
	.Selector4(\hps_0_h2f_axi_master_agent|Selector4~1_combout ),
	.Add3(\hps_0_h2f_axi_master_agent|Add3~1_combout ),
	.Add31(\hps_0_h2f_axi_master_agent|Add3~2_combout ),
	.Selector11(\hps_0_h2f_axi_master_agent|Selector11~0_combout ),
	.Selector111(\hps_0_h2f_axi_master_agent|Selector11~1_combout ),
	.base_address_2(\hps_0_h2f_axi_master_agent|align_address_to_size|base_address[2]~1_combout ),
	.Selector5(\hps_0_h2f_axi_master_agent|Selector5~1_combout ),
	.Add32(\hps_0_h2f_axi_master_agent|Add3~3_combout ),
	.Selector12(\hps_0_h2f_axi_master_agent|Selector12~0_combout ),
	.out_data_1(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[1]~5_combout ),
	.out_data_0(\hps_0_h2f_axi_master_agent|align_address_to_size|out_data[0]~6_combout ),
	.Selector6(\hps_0_h2f_axi_master_agent|Selector6~0_combout ),
	.Selector13(\hps_0_h2f_axi_master_agent|Selector13~1_combout ),
	.clk_clk(clk_clk));

spw_babasu_altera_merlin_slave_translator_9 spill_enable_s1_translator(
	.waitrequest_reset_override(\autostart_s1_translator|waitrequest_reset_override~q ),
	.out_valid_reg(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\spill_enable_s1_agent_rsp_fifo|mem_used[1]~q ),
	.WideOr0(\spill_enable_s1_agent|WideOr0~0_combout ),
	.wait_latency_counter_1(wait_latency_counter_12),
	.wait_latency_counter_0(wait_latency_counter_02),
	.read_latency_shift_reg_0(\spill_enable_s1_translator|read_latency_shift_reg[0]~q ),
	.av_readdata_pre_0(\spill_enable_s1_translator|av_readdata_pre[0]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.m0_write(m0_write5),
	.cp_ready(\spill_enable_s1_agent|cp_ready~3_combout ),
	.in_data_reg_69(\spill_enable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_014}),
	.clk(clk_clk));

spw_babasu_altera_merlin_slave_translator_14 tx_clk_div_s1_translator(
	.waitrequest_reset_override(\autostart_s1_translator|waitrequest_reset_override~q ),
	.out_valid_reg(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\tx_clk_div_s1_agent_rsp_fifo|mem_used[1]~q ),
	.WideOr0(\tx_clk_div_s1_agent|WideOr0~0_combout ),
	.wait_latency_counter_1(wait_latency_counter_11),
	.wait_latency_counter_0(wait_latency_counter_01),
	.read_latency_shift_reg_0(\tx_clk_div_s1_translator|read_latency_shift_reg[0]~q ),
	.av_readdata_pre_0(\tx_clk_div_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\tx_clk_div_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\tx_clk_div_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\tx_clk_div_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\tx_clk_div_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\tx_clk_div_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_6(\tx_clk_div_s1_translator|av_readdata_pre[6]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.m0_write(m0_write8),
	.cp_ready(\tx_clk_div_s1_agent|cp_ready~4_combout ),
	.in_data_reg_69(\tx_clk_div_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_65,readdata_55,readdata_45,readdata_35,readdata_26,readdata_16,readdata_01}),
	.clk(clk_clk));

spw_babasu_altera_merlin_slave_translator_12 time_in_s1_translator(
	.waitrequest_reset_override(\autostart_s1_translator|waitrequest_reset_override~q ),
	.out_valid_reg(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\time_in_s1_agent_rsp_fifo|mem_used[1]~q ),
	.WideOr0(\time_in_s1_agent|WideOr0~0_combout ),
	.wait_latency_counter_1(wait_latency_counter_14),
	.wait_latency_counter_0(wait_latency_counter_04),
	.read_latency_shift_reg_0(\time_in_s1_translator|read_latency_shift_reg[0]~q ),
	.av_readdata_pre_0(\time_in_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\time_in_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\time_in_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\time_in_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\time_in_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\time_in_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_6(\time_in_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_7(\time_in_s1_translator|av_readdata_pre[7]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.m0_write(m0_write7),
	.cp_ready(\time_in_s1_agent|cp_ready~4_combout ),
	.in_data_reg_69(\time_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_72,readdata_64,readdata_54,readdata_44,readdata_34,readdata_25,readdata_15,readdata_016}),
	.clk(clk_clk));

spw_babasu_altera_merlin_slave_translator_10 tick_in_s1_translator(
	.waitrequest_reset_override(\autostart_s1_translator|waitrequest_reset_override~q ),
	.out_valid_reg(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\tick_in_s1_agent_rsp_fifo|mem_used[1]~q ),
	.WideOr0(\tick_in_s1_agent|WideOr0~0_combout ),
	.wait_latency_counter_1(wait_latency_counter_13),
	.wait_latency_counter_0(wait_latency_counter_03),
	.read_latency_shift_reg_0(\tick_in_s1_translator|read_latency_shift_reg[0]~q ),
	.av_readdata_pre_0(\tick_in_s1_translator|av_readdata_pre[0]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.m0_write(m0_write6),
	.cp_ready(\tick_in_s1_agent|cp_ready~4_combout ),
	.in_data_reg_69(\tick_in_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_013}),
	.clk(clk_clk));

spw_babasu_altera_merlin_slave_translator_13 time_out_s1_translator(
	.wait_latency_counter_1(\time_out_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\time_out_s1_translator|wait_latency_counter[0]~q ),
	.read_latency_shift_reg_0(\time_out_s1_translator|read_latency_shift_reg[0]~q ),
	.av_readdata_pre_0(\time_out_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\time_out_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\time_out_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\time_out_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\time_out_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\time_out_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_6(\time_out_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_7(\time_out_s1_translator|av_readdata_pre[7]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.write(\time_out_s1_agent_rsp_fifo|write~0_combout ),
	.write1(\time_out_s1_agent_rsp_fifo|write~1_combout ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_73,readdata_62,readdata_52,readdata_42,readdata_32,readdata_22,readdata_12,readdata_06}),
	.clk(clk_clk));

spw_babasu_altera_merlin_slave_translator_11 tick_out_s1_translator(
	.wait_latency_counter_1(\tick_out_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\tick_out_s1_translator|wait_latency_counter[0]~q ),
	.read_latency_shift_reg_0(\tick_out_s1_translator|read_latency_shift_reg[0]~q ),
	.av_readdata_pre_0(\tick_out_s1_translator|av_readdata_pre[0]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.write(\tick_out_s1_agent_rsp_fifo|write~0_combout ),
	.write1(\tick_out_s1_agent_rsp_fifo|write~1_combout ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_07}),
	.clk(clk_clk));

spw_babasu_altera_merlin_slave_translator_8 rx_empty_s1_translator(
	.wait_latency_counter_1(\rx_empty_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\rx_empty_s1_translator|wait_latency_counter[0]~q ),
	.read_latency_shift_reg_0(\rx_empty_s1_translator|read_latency_shift_reg[0]~q ),
	.av_readdata_pre_0(\rx_empty_s1_translator|av_readdata_pre[0]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.write(\rx_empty_s1_agent_rsp_fifo|write~0_combout ),
	.write1(\rx_empty_s1_agent_rsp_fifo|write~1_combout ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_08}),
	.clk(clk_clk));

spw_babasu_altera_merlin_slave_translator_6 link_start_s1_translator(
	.waitrequest_reset_override(\autostart_s1_translator|waitrequest_reset_override~q ),
	.out_valid_reg(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\link_start_s1_agent_rsp_fifo|mem_used[1]~q ),
	.WideOr0(\link_start_s1_agent|WideOr0~0_combout ),
	.wait_latency_counter_1(wait_latency_counter_17),
	.wait_latency_counter_0(wait_latency_counter_07),
	.read_latency_shift_reg_0(\link_start_s1_translator|read_latency_shift_reg[0]~q ),
	.av_readdata_pre_0(\link_start_s1_translator|av_readdata_pre[0]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.m0_write(m0_write3),
	.cp_ready(\link_start_s1_agent|cp_ready~3_combout ),
	.in_data_reg_69(\link_start_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_09}),
	.clk(clk_clk));

spw_babasu_altera_merlin_slave_translator_7 rd_data_s1_translator(
	.waitrequest_reset_override(\autostart_s1_translator|waitrequest_reset_override~q ),
	.out_valid_reg(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\rd_data_s1_agent_rsp_fifo|mem_used[1]~q ),
	.WideOr0(\rd_data_s1_agent|WideOr0~0_combout ),
	.wait_latency_counter_1(wait_latency_counter_16),
	.wait_latency_counter_0(wait_latency_counter_06),
	.read_latency_shift_reg_0(\rd_data_s1_translator|read_latency_shift_reg[0]~q ),
	.av_readdata_pre_0(\rd_data_s1_translator|av_readdata_pre[0]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.m0_write(m0_write4),
	.cp_ready(\rd_data_s1_agent|cp_ready~4_combout ),
	.in_data_reg_69(\rd_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_012}),
	.clk(clk_clk));

spw_babasu_altera_merlin_slave_translator_3 data_o_s1_translator(
	.wait_latency_counter_1(\data_o_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\data_o_s1_translator|wait_latency_counter[0]~q ),
	.read_latency_shift_reg_0(\data_o_s1_translator|read_latency_shift_reg[0]~q ),
	.av_readdata_pre_0(\data_o_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\data_o_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\data_o_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\data_o_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\data_o_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\data_o_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_6(\data_o_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_7(\data_o_s1_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_8(\data_o_s1_translator|av_readdata_pre[8]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.write(\data_o_s1_agent_rsp_fifo|write~0_combout ),
	.write1(\data_o_s1_agent_rsp_fifo|write~1_combout ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_82,readdata_74,readdata_63,readdata_53,readdata_43,readdata_33,readdata_23,readdata_13,readdata_03}),
	.clk(clk_clk));

spw_babasu_altera_merlin_slave_translator_15 tx_full_s1_translator(
	.wait_latency_counter_1(\tx_full_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\tx_full_s1_translator|wait_latency_counter[0]~q ),
	.read_latency_shift_reg_0(\tx_full_s1_translator|read_latency_shift_reg[0]~q ),
	.av_readdata_pre_0(\tx_full_s1_translator|av_readdata_pre[0]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.write(\tx_full_s1_agent_rsp_fifo|write~0_combout ),
	.write1(\tx_full_s1_agent_rsp_fifo|write~1_combout ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_04}),
	.clk(clk_clk));

spw_babasu_altera_merlin_slave_translator_16 wr_data_s1_translator(
	.waitrequest_reset_override(\autostart_s1_translator|waitrequest_reset_override~q ),
	.out_valid_reg(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\wr_data_s1_agent_rsp_fifo|mem_used[1]~q ),
	.WideOr0(\wr_data_s1_agent|WideOr0~0_combout ),
	.wait_latency_counter_1(wait_latency_counter_19),
	.wait_latency_counter_0(wait_latency_counter_09),
	.read_latency_shift_reg_0(\wr_data_s1_translator|read_latency_shift_reg[0]~q ),
	.av_readdata_pre_0(\wr_data_s1_translator|av_readdata_pre[0]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.m0_write(m0_write9),
	.cp_ready(\wr_data_s1_agent|cp_ready~4_combout ),
	.in_data_reg_69(\wr_data_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_011}),
	.clk(clk_clk));

spw_babasu_altera_merlin_slave_translator_2 data_i_s1_translator(
	.waitrequest_reset_override(\autostart_s1_translator|waitrequest_reset_override~q ),
	.out_valid_reg(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\data_i_s1_agent_rsp_fifo|mem_used[1]~q ),
	.WideOr0(\data_i_s1_agent|WideOr0~0_combout ),
	.wait_latency_counter_1(wait_latency_counter_15),
	.wait_latency_counter_0(wait_latency_counter_05),
	.read_latency_shift_reg_0(\data_i_s1_translator|read_latency_shift_reg[0]~q ),
	.av_readdata_pre_0(\data_i_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\data_i_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\data_i_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\data_i_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\data_i_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\data_i_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_6(\data_i_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_7(\data_i_s1_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_8(\data_i_s1_translator|av_readdata_pre[8]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.m0_write(m0_write1),
	.cp_ready(\data_i_s1_agent|cp_ready~4_combout ),
	.in_data_reg_69(\data_i_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_8,readdata_71,readdata_61,readdata_51,readdata_41,readdata_31,readdata_21,readdata_11,readdata_015}),
	.clk(clk_clk));

spw_babasu_altera_merlin_slave_translator_4 flags_s1_translator(
	.wait_latency_counter_1(\flags_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\flags_s1_translator|wait_latency_counter[0]~q ),
	.read_latency_shift_reg_0(\flags_s1_translator|read_latency_shift_reg[0]~q ),
	.av_readdata_pre_0(\flags_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\flags_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\flags_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\flags_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\flags_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\flags_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_6(\flags_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_7(\flags_s1_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_8(\flags_s1_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_9(\flags_s1_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_10(\flags_s1_translator|av_readdata_pre[10]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.write(\flags_s1_agent_rsp_fifo|write~0_combout ),
	.write1(\flags_s1_agent_rsp_fifo|write~1_combout ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_10,readdata_9,readdata_81,readdata_7,readdata_6,readdata_5,readdata_4,readdata_3,readdata_24,readdata_14,readdata_05}),
	.clk(clk_clk));

spw_babasu_altera_merlin_slave_translator_1 currentstate_s1_translator(
	.wait_latency_counter_1(\currentstate_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\currentstate_s1_translator|wait_latency_counter[0]~q ),
	.read_latency_shift_reg_0(\currentstate_s1_translator|read_latency_shift_reg[0]~q ),
	.av_readdata_pre_0(\currentstate_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\currentstate_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\currentstate_s1_translator|av_readdata_pre[2]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.write(\currentstate_s1_agent_rsp_fifo|write~0_combout ),
	.write1(\currentstate_s1_agent_rsp_fifo|write~1_combout ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_2,readdata_1,readdata_02}),
	.clk(clk_clk));

spw_babasu_altera_merlin_slave_translator autostart_s1_translator(
	.waitrequest_reset_override1(\autostart_s1_translator|waitrequest_reset_override~q ),
	.out_valid_reg(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\autostart_s1_agent_rsp_fifo|mem_used[1]~q ),
	.WideOr0(\autostart_s1_agent|WideOr0~0_combout ),
	.wait_latency_counter_1(wait_latency_counter_18),
	.wait_latency_counter_0(wait_latency_counter_08),
	.read_latency_shift_reg_0(\autostart_s1_translator|read_latency_shift_reg[0]~q ),
	.av_readdata_pre_0(\autostart_s1_translator|av_readdata_pre[0]~q ),
	.m0_write(m0_write),
	.reset(altera_reset_synchronizer_int_chain_out),
	.cp_ready(\autostart_s1_agent|cp_ready~4_combout ),
	.in_data_reg_69(\autostart_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_0}),
	.clk(clk_clk));

spw_babasu_altera_merlin_slave_translator_5 link_disable_s1_translator(
	.waitrequest_reset_override(\autostart_s1_translator|waitrequest_reset_override~q ),
	.out_valid_reg(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\link_disable_s1_agent_rsp_fifo|mem_used[1]~q ),
	.WideOr0(\link_disable_s1_agent|WideOr0~0_combout ),
	.wait_latency_counter_1(wait_latency_counter_1),
	.wait_latency_counter_0(wait_latency_counter_0),
	.read_latency_shift_reg_0(\link_disable_s1_translator|read_latency_shift_reg[0]~q ),
	.av_readdata_pre_0(\link_disable_s1_translator|av_readdata_pre[0]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.m0_write(m0_write2),
	.cp_ready(\link_disable_s1_agent|cp_ready~4_combout ),
	.in_data_reg_69(\link_disable_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_010}),
	.clk(clk_clk));

endmodule

module spw_babasu_altera_avalon_sc_fifo (
	read_latency_shift_reg_0,
	mem_used_0,
	mem_129_0,
	mem_used_01,
	av_readdata_pre_0,
	mem_0_0,
	reset,
	WideOr0,
	clk)/* synthesis synthesis_greybox=0 */;
input 	read_latency_shift_reg_0;
output 	mem_used_0;
input 	mem_129_0;
input 	mem_used_01;
input 	av_readdata_pre_0;
output 	mem_0_0;
input 	reset;
input 	WideOr0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~q ;
wire \mem_used[0]~0_combout ;
wire \mem[1][0]~q ;
wire \mem~0_combout ;
wire \mem[0][0]~1_combout ;


dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][0] (
	.clk(clk),
	.d(\mem[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_0_0),
	.prn(vcc));
defparam \mem[0][0] .is_wysiwyg = "true";
defparam \mem[0][0] .power_up = "low";

cyclonev_lcell_comb \read~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_129_0),
	.datad(!mem_used_01),
	.datae(!WideOr0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h0000777000007770;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!\mem_used[1]~q ),
	.datad(!\read~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'h1F001F001F001F00;
defparam \mem_used[1]~1 .shared_arith = "off";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[1]~q ),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!\mem_used[1]~q ),
	.datad(!\read~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~0 .extended_lut = "off";
defparam \mem_used[0]~0 .lut_mask = 64'h731F731F731F731F;
defparam \mem_used[0]~0 .shared_arith = "off";

dffeas \mem[1][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][0]~q ),
	.prn(vcc));
defparam \mem[1][0] .is_wysiwyg = "true";
defparam \mem[1][0] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!av_readdata_pre_0),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h4747474747474747;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \mem[0][0]~1 (
	.dataa(!mem_used_0),
	.datab(!mem_0_0),
	.datac(!\read~0_combout ),
	.datad(!\mem~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem[0][0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem[0][0]~1 .extended_lut = "off";
defparam \mem[0][0]~1 .lut_mask = 64'h10BF10BF10BF10BF;
defparam \mem[0][0]~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_avalon_sc_fifo_1 (
	out_valid_reg,
	mem_used_1,
	WideOr0,
	in_data_reg_68,
	stateST_UNCOMP_WR_SUBBURST,
	mem_129_0,
	mem_used_0,
	mem_68_0,
	mem_66_0,
	comb,
	mem_130_0,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	mem_105_0,
	mem_106_0,
	mem_107_0,
	mem_108_0,
	mem_109_0,
	mem_110_0,
	mem_111_0,
	mem_112_0,
	mem_113_0,
	mem_114_0,
	mem_115_0,
	mem_116_0,
	reset,
	nxt_out_eop,
	last_packet_beat,
	WideOr01,
	read,
	cp_ready,
	in_data_reg_69,
	rf_source_valid,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_6,
	sink_ready,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	clk)/* synthesis synthesis_greybox=0 */;
input 	out_valid_reg;
output 	mem_used_1;
input 	WideOr0;
input 	in_data_reg_68;
input 	stateST_UNCOMP_WR_SUBBURST;
output 	mem_129_0;
output 	mem_used_0;
output 	mem_68_0;
output 	mem_66_0;
input 	comb;
output 	mem_130_0;
output 	mem_78_0;
output 	mem_77_0;
output 	mem_76_0;
output 	mem_75_0;
output 	mem_74_0;
output 	mem_105_0;
output 	mem_106_0;
output 	mem_107_0;
output 	mem_108_0;
output 	mem_109_0;
output 	mem_110_0;
output 	mem_111_0;
output 	mem_112_0;
output 	mem_113_0;
output 	mem_114_0;
output 	mem_115_0;
output 	mem_116_0;
input 	reset;
input 	nxt_out_eop;
input 	last_packet_beat;
input 	WideOr01;
output 	read;
input 	cp_ready;
input 	in_data_reg_69;
input 	rf_source_valid;
input 	out_byte_cnt_reg_2;
input 	out_uncomp_byte_cnt_reg_5;
input 	out_uncomp_byte_cnt_reg_4;
input 	out_uncomp_byte_cnt_reg_3;
input 	out_uncomp_byte_cnt_reg_2;
input 	out_uncomp_byte_cnt_reg_6;
input 	sink_ready;
input 	in_data_reg_105;
input 	in_data_reg_106;
input 	in_data_reg_107;
input 	in_data_reg_108;
input 	in_data_reg_109;
input 	in_data_reg_110;
input 	in_data_reg_111;
input 	in_data_reg_112;
input 	in_data_reg_113;
input 	in_data_reg_114;
input 	in_data_reg_115;
input 	in_data_reg_116;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \write~0_combout ;
wire \mem_used[1]~0_combout ;
wire \mem[1][129]~q ;
wire \mem~20_combout ;
wire \always0~0_combout ;
wire \mem_used[0]~1_combout ;
wire \mem[1][68]~q ;
wire \mem~0_combout ;
wire \mem[1][69]~q ;
wire \mem~1_combout ;
wire \mem[1][130]~q ;
wire \mem~2_combout ;
wire \mem[1][78]~q ;
wire \mem~3_combout ;
wire \mem[1][77]~q ;
wire \mem~4_combout ;
wire \mem[1][76]~q ;
wire \mem~5_combout ;
wire \mem[1][75]~q ;
wire \mem~6_combout ;
wire \mem[1][74]~q ;
wire \mem~7_combout ;
wire \mem[1][105]~q ;
wire \mem~8_combout ;
wire \mem[1][106]~q ;
wire \mem~9_combout ;
wire \mem[1][107]~q ;
wire \mem~10_combout ;
wire \mem[1][108]~q ;
wire \mem~11_combout ;
wire \mem[1][109]~q ;
wire \mem~12_combout ;
wire \mem[1][110]~q ;
wire \mem~13_combout ;
wire \mem[1][111]~q ;
wire \mem~14_combout ;
wire \mem[1][112]~q ;
wire \mem~15_combout ;
wire \mem[1][113]~q ;
wire \mem~16_combout ;
wire \mem[1][114]~q ;
wire \mem~17_combout ;
wire \mem[1][115]~q ;
wire \mem~18_combout ;
wire \mem[1][116]~q ;
wire \mem~19_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][129] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_129_0),
	.prn(vcc));
defparam \mem[0][129] .is_wysiwyg = "true";
defparam \mem[0][129] .power_up = "low";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][68] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_68_0),
	.prn(vcc));
defparam \mem[0][68] .is_wysiwyg = "true";
defparam \mem[0][68] .power_up = "low";

dffeas \mem[0][66] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_66_0),
	.prn(vcc));
defparam \mem[0][66] .is_wysiwyg = "true";
defparam \mem[0][66] .power_up = "low";

dffeas \mem[0][130] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_130_0),
	.prn(vcc));
defparam \mem[0][130] .is_wysiwyg = "true";
defparam \mem[0][130] .power_up = "low";

dffeas \mem[0][78] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_78_0),
	.prn(vcc));
defparam \mem[0][78] .is_wysiwyg = "true";
defparam \mem[0][78] .power_up = "low";

dffeas \mem[0][77] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_77_0),
	.prn(vcc));
defparam \mem[0][77] .is_wysiwyg = "true";
defparam \mem[0][77] .power_up = "low";

dffeas \mem[0][76] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_76_0),
	.prn(vcc));
defparam \mem[0][76] .is_wysiwyg = "true";
defparam \mem[0][76] .power_up = "low";

dffeas \mem[0][75] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_75_0),
	.prn(vcc));
defparam \mem[0][75] .is_wysiwyg = "true";
defparam \mem[0][75] .power_up = "low";

dffeas \mem[0][74] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_74_0),
	.prn(vcc));
defparam \mem[0][74] .is_wysiwyg = "true";
defparam \mem[0][74] .power_up = "low";

dffeas \mem[0][105] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_105_0),
	.prn(vcc));
defparam \mem[0][105] .is_wysiwyg = "true";
defparam \mem[0][105] .power_up = "low";

dffeas \mem[0][106] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_106_0),
	.prn(vcc));
defparam \mem[0][106] .is_wysiwyg = "true";
defparam \mem[0][106] .power_up = "low";

dffeas \mem[0][107] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_107_0),
	.prn(vcc));
defparam \mem[0][107] .is_wysiwyg = "true";
defparam \mem[0][107] .power_up = "low";

dffeas \mem[0][108] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_108_0),
	.prn(vcc));
defparam \mem[0][108] .is_wysiwyg = "true";
defparam \mem[0][108] .power_up = "low";

dffeas \mem[0][109] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_109_0),
	.prn(vcc));
defparam \mem[0][109] .is_wysiwyg = "true";
defparam \mem[0][109] .power_up = "low";

dffeas \mem[0][110] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_110_0),
	.prn(vcc));
defparam \mem[0][110] .is_wysiwyg = "true";
defparam \mem[0][110] .power_up = "low";

dffeas \mem[0][111] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_111_0),
	.prn(vcc));
defparam \mem[0][111] .is_wysiwyg = "true";
defparam \mem[0][111] .power_up = "low";

dffeas \mem[0][112] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_112_0),
	.prn(vcc));
defparam \mem[0][112] .is_wysiwyg = "true";
defparam \mem[0][112] .power_up = "low";

dffeas \mem[0][113] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_113_0),
	.prn(vcc));
defparam \mem[0][113] .is_wysiwyg = "true";
defparam \mem[0][113] .power_up = "low";

dffeas \mem[0][114] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_114_0),
	.prn(vcc));
defparam \mem[0][114] .is_wysiwyg = "true";
defparam \mem[0][114] .power_up = "low";

dffeas \mem[0][115] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_115_0),
	.prn(vcc));
defparam \mem[0][115] .is_wysiwyg = "true";
defparam \mem[0][115] .power_up = "low";

dffeas \mem[0][116] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_116_0),
	.prn(vcc));
defparam \mem[0][116] .is_wysiwyg = "true";
defparam \mem[0][116] .power_up = "low";

cyclonev_lcell_comb \read~0 (
	.dataa(!comb),
	.datab(!WideOr01),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h1111111111111111;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \write~0 (
	.dataa(!mem_used_1),
	.datab(!WideOr0),
	.datac(!cp_ready),
	.datad(!rf_source_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'h008A008A008A008A;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!last_packet_beat),
	.datad(!read),
	.datae(!\write~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'h5505335355053353;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][129] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][129]~q ),
	.prn(vcc));
defparam \mem[1][129] .is_wysiwyg = "true";
defparam \mem[1][129] .power_up = "low";

cyclonev_lcell_comb \mem~20 (
	.dataa(!WideOr0),
	.datab(!out_valid_reg),
	.datac(!\mem[1][129]~q ),
	.datad(!in_data_reg_68),
	.datae(!mem_used_1),
	.dataf(!nxt_out_eop),
	.datag(!in_data_reg_69),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~20 .extended_lut = "on";
defparam \mem~20 .lut_mask = 64'h02020F0F02330F0F;
defparam \mem~20 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!mem_used_0),
	.datab(!sink_ready),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!\write~0_combout ),
	.datad(!sink_ready),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'h3F1F3F1F3F1F3F1F;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem[1][68] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][68]~q ),
	.prn(vcc));
defparam \mem[1][68] .is_wysiwyg = "true";
defparam \mem[1][68] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!mem_used_1),
	.datab(!in_data_reg_68),
	.datac(!\mem[1][68]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h2727272727272727;
defparam \mem~0 .shared_arith = "off";

dffeas \mem[1][69] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][69]~q ),
	.prn(vcc));
defparam \mem[1][69] .is_wysiwyg = "true";
defparam \mem[1][69] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!mem_used_1),
	.datab(!in_data_reg_69),
	.datac(!\mem[1][69]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h2727272727272727;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[1][130] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][130]~q ),
	.prn(vcc));
defparam \mem[1][130] .is_wysiwyg = "true";
defparam \mem[1][130] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!mem_used_1),
	.datab(!nxt_out_eop),
	.datac(!\mem[1][130]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h2727272727272727;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[1][78] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][78]~q ),
	.prn(vcc));
defparam \mem[1][78] .is_wysiwyg = "true";
defparam \mem[1][78] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_6),
	.datad(!\mem[1][78]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h0257025702570257;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][77] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][77]~q ),
	.prn(vcc));
defparam \mem[1][77] .is_wysiwyg = "true";
defparam \mem[1][77] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\mem[1][77]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h0257025702570257;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][76] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][76]~q ),
	.prn(vcc));
defparam \mem[1][76] .is_wysiwyg = "true";
defparam \mem[1][76] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!\mem[1][76]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h0257025702570257;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][75] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][75]~q ),
	.prn(vcc));
defparam \mem[1][75] .is_wysiwyg = "true";
defparam \mem[1][75] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\mem[1][75]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h0257025702570257;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[1][74] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][74]~q ),
	.prn(vcc));
defparam \mem[1][74] .is_wysiwyg = "true";
defparam \mem[1][74] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_byte_cnt_reg_2),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(!\mem[1][74]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h082A5D7F082A5D7F;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[1][105] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][105]~q ),
	.prn(vcc));
defparam \mem[1][105] .is_wysiwyg = "true";
defparam \mem[1][105] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][105]~q ),
	.datac(!in_data_reg_105),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~8 .shared_arith = "off";

dffeas \mem[1][106] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][106]~q ),
	.prn(vcc));
defparam \mem[1][106] .is_wysiwyg = "true";
defparam \mem[1][106] .power_up = "low";

cyclonev_lcell_comb \mem~9 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][106]~q ),
	.datac(!in_data_reg_106),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~9 .extended_lut = "off";
defparam \mem~9 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~9 .shared_arith = "off";

dffeas \mem[1][107] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][107]~q ),
	.prn(vcc));
defparam \mem[1][107] .is_wysiwyg = "true";
defparam \mem[1][107] .power_up = "low";

cyclonev_lcell_comb \mem~10 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][107]~q ),
	.datac(!in_data_reg_107),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~10 .extended_lut = "off";
defparam \mem~10 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~10 .shared_arith = "off";

dffeas \mem[1][108] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][108]~q ),
	.prn(vcc));
defparam \mem[1][108] .is_wysiwyg = "true";
defparam \mem[1][108] .power_up = "low";

cyclonev_lcell_comb \mem~11 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][108]~q ),
	.datac(!in_data_reg_108),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~11 .extended_lut = "off";
defparam \mem~11 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~11 .shared_arith = "off";

dffeas \mem[1][109] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][109]~q ),
	.prn(vcc));
defparam \mem[1][109] .is_wysiwyg = "true";
defparam \mem[1][109] .power_up = "low";

cyclonev_lcell_comb \mem~12 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][109]~q ),
	.datac(!in_data_reg_109),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~12 .extended_lut = "off";
defparam \mem~12 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~12 .shared_arith = "off";

dffeas \mem[1][110] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][110]~q ),
	.prn(vcc));
defparam \mem[1][110] .is_wysiwyg = "true";
defparam \mem[1][110] .power_up = "low";

cyclonev_lcell_comb \mem~13 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][110]~q ),
	.datac(!in_data_reg_110),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~13 .extended_lut = "off";
defparam \mem~13 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~13 .shared_arith = "off";

dffeas \mem[1][111] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][111]~q ),
	.prn(vcc));
defparam \mem[1][111] .is_wysiwyg = "true";
defparam \mem[1][111] .power_up = "low";

cyclonev_lcell_comb \mem~14 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][111]~q ),
	.datac(!in_data_reg_111),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~14 .extended_lut = "off";
defparam \mem~14 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~14 .shared_arith = "off";

dffeas \mem[1][112] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][112]~q ),
	.prn(vcc));
defparam \mem[1][112] .is_wysiwyg = "true";
defparam \mem[1][112] .power_up = "low";

cyclonev_lcell_comb \mem~15 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][112]~q ),
	.datac(!in_data_reg_112),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~15 .extended_lut = "off";
defparam \mem~15 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~15 .shared_arith = "off";

dffeas \mem[1][113] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][113]~q ),
	.prn(vcc));
defparam \mem[1][113] .is_wysiwyg = "true";
defparam \mem[1][113] .power_up = "low";

cyclonev_lcell_comb \mem~16 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][113]~q ),
	.datac(!in_data_reg_113),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~16 .extended_lut = "off";
defparam \mem~16 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~16 .shared_arith = "off";

dffeas \mem[1][114] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][114]~q ),
	.prn(vcc));
defparam \mem[1][114] .is_wysiwyg = "true";
defparam \mem[1][114] .power_up = "low";

cyclonev_lcell_comb \mem~17 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][114]~q ),
	.datac(!in_data_reg_114),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~17 .extended_lut = "off";
defparam \mem~17 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~17 .shared_arith = "off";

dffeas \mem[1][115] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][115]~q ),
	.prn(vcc));
defparam \mem[1][115] .is_wysiwyg = "true";
defparam \mem[1][115] .power_up = "low";

cyclonev_lcell_comb \mem~18 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][115]~q ),
	.datac(!in_data_reg_115),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~18 .extended_lut = "off";
defparam \mem~18 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~18 .shared_arith = "off";

dffeas \mem[1][116] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][116]~q ),
	.prn(vcc));
defparam \mem[1][116] .is_wysiwyg = "true";
defparam \mem[1][116] .power_up = "low";

cyclonev_lcell_comb \mem~19 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][116]~q ),
	.datac(!in_data_reg_116),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~19 .extended_lut = "off";
defparam \mem~19 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~19 .shared_arith = "off";

endmodule

module spw_babasu_altera_avalon_sc_fifo_2 (
	h2f_RREADY_0,
	read_latency_shift_reg_0,
	mem_used_0,
	empty1,
	av_readdata_pre_0,
	mem_0_0,
	av_readdata_pre_1,
	mem_1_0,
	av_readdata_pre_2,
	mem_2_0,
	reset,
	clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_RREADY_0;
input 	read_latency_shift_reg_0;
output 	mem_used_0;
output 	empty1;
input 	av_readdata_pre_0;
output 	mem_0_0;
input 	av_readdata_pre_1;
output 	mem_1_0;
input 	av_readdata_pre_2;
output 	mem_2_0;
input 	reset;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[1]~1_combout ;
wire \mem_used[1]~q ;
wire \mem_used[0]~0_combout ;
wire \mem[1][0]~q ;
wire \mem~0_combout ;
wire \always0~0_combout ;
wire \mem[1][1]~q ;
wire \mem~1_combout ;
wire \mem[1][2]~q ;
wire \mem~2_combout ;


dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb empty(
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(empty1),
	.sumout(),
	.cout(),
	.shareout());
defparam empty.extended_lut = "off";
defparam empty.lut_mask = 64'h8888888888888888;
defparam empty.shared_arith = "off";

dffeas \mem[0][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_0_0),
	.prn(vcc));
defparam \mem[0][0] .is_wysiwyg = "true";
defparam \mem[0][0] .power_up = "low";

dffeas \mem[0][1] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_1_0),
	.prn(vcc));
defparam \mem[0][1] .is_wysiwyg = "true";
defparam \mem[0][1] .power_up = "low";

dffeas \mem[0][2] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_2_0),
	.prn(vcc));
defparam \mem[0][2] .is_wysiwyg = "true";
defparam \mem[0][2] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!h2f_RREADY_0),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem_used[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'h02EA02EA02EA02EA;
defparam \mem_used[1]~1 .shared_arith = "off";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[1]~q ),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~0 (
	.dataa(!h2f_RREADY_0),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem_used[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~0 .extended_lut = "off";
defparam \mem_used[0]~0 .lut_mask = 64'h2B1F2B1F2B1F2B1F;
defparam \mem_used[0]~0 .shared_arith = "off";

dffeas \mem[1][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][0]~q ),
	.prn(vcc));
defparam \mem[1][0] .is_wysiwyg = "true";
defparam \mem[1][0] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!av_readdata_pre_0),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h4747474747474747;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!h2f_RREADY_0),
	.datab(!mem_used_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \always0~0 .shared_arith = "off";

dffeas \mem[1][1] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][1]~q ),
	.prn(vcc));
defparam \mem[1][1] .is_wysiwyg = "true";
defparam \mem[1][1] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!av_readdata_pre_1),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h4747474747474747;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[1][2] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][2]~q ),
	.prn(vcc));
defparam \mem[1][2] .is_wysiwyg = "true";
defparam \mem[1][2] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!av_readdata_pre_2),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h4747474747474747;
defparam \mem~2 .shared_arith = "off";

endmodule

module spw_babasu_altera_avalon_sc_fifo_3 (
	h2f_RREADY_0,
	waitrequest_reset_override,
	mem_used_1,
	in_data_reg_69,
	wait_latency_counter_1,
	wait_latency_counter_0,
	nxt_out_eop,
	out_valid_reg,
	stateST_UNCOMP_WR_SUBBURST,
	mem_130_0,
	empty,
	mem_66_0,
	mem_used_0,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	mem_105_0,
	mem_106_0,
	mem_107_0,
	mem_108_0,
	mem_109_0,
	mem_110_0,
	mem_111_0,
	mem_112_0,
	mem_113_0,
	mem_114_0,
	mem_115_0,
	mem_116_0,
	reset,
	last_packet_beat,
	write,
	write1,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_6,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_RREADY_0;
input 	waitrequest_reset_override;
output 	mem_used_1;
input 	in_data_reg_69;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	nxt_out_eop;
input 	out_valid_reg;
input 	stateST_UNCOMP_WR_SUBBURST;
output 	mem_130_0;
input 	empty;
output 	mem_66_0;
output 	mem_used_0;
output 	mem_78_0;
output 	mem_77_0;
output 	mem_76_0;
output 	mem_75_0;
output 	mem_74_0;
output 	mem_105_0;
output 	mem_106_0;
output 	mem_107_0;
output 	mem_108_0;
output 	mem_109_0;
output 	mem_110_0;
output 	mem_111_0;
output 	mem_112_0;
output 	mem_113_0;
output 	mem_114_0;
output 	mem_115_0;
output 	mem_116_0;
input 	reset;
input 	last_packet_beat;
output 	write;
output 	write1;
input 	out_byte_cnt_reg_2;
input 	out_uncomp_byte_cnt_reg_3;
input 	out_uncomp_byte_cnt_reg_2;
input 	out_uncomp_byte_cnt_reg_4;
input 	out_uncomp_byte_cnt_reg_5;
input 	out_uncomp_byte_cnt_reg_6;
input 	in_data_reg_105;
input 	in_data_reg_106;
input 	in_data_reg_107;
input 	in_data_reg_108;
input 	in_data_reg_109;
input 	in_data_reg_110;
input 	in_data_reg_111;
input 	in_data_reg_112;
input 	in_data_reg_113;
input 	in_data_reg_114;
input 	in_data_reg_115;
input 	in_data_reg_116;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read~0_combout ;
wire \mem_used[1]~0_combout ;
wire \mem[1][130]~q ;
wire \mem~0_combout ;
wire \always0~0_combout ;
wire \mem[1][69]~q ;
wire \mem~1_combout ;
wire \mem_used[0]~1_combout ;
wire \mem[1][78]~q ;
wire \mem~2_combout ;
wire \mem[1][77]~q ;
wire \mem~3_combout ;
wire \mem[1][76]~q ;
wire \mem~4_combout ;
wire \mem[1][75]~q ;
wire \mem~5_combout ;
wire \mem[1][74]~q ;
wire \mem~6_combout ;
wire \mem[1][105]~q ;
wire \mem~7_combout ;
wire \mem[1][106]~q ;
wire \mem~8_combout ;
wire \mem[1][107]~q ;
wire \mem~9_combout ;
wire \mem[1][108]~q ;
wire \mem~10_combout ;
wire \mem[1][109]~q ;
wire \mem~11_combout ;
wire \mem[1][110]~q ;
wire \mem~12_combout ;
wire \mem[1][111]~q ;
wire \mem~13_combout ;
wire \mem[1][112]~q ;
wire \mem~14_combout ;
wire \mem[1][113]~q ;
wire \mem~15_combout ;
wire \mem[1][114]~q ;
wire \mem~16_combout ;
wire \mem[1][115]~q ;
wire \mem~17_combout ;
wire \mem[1][116]~q ;
wire \mem~18_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][130] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_130_0),
	.prn(vcc));
defparam \mem[0][130] .is_wysiwyg = "true";
defparam \mem[0][130] .power_up = "low";

dffeas \mem[0][66] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_66_0),
	.prn(vcc));
defparam \mem[0][66] .is_wysiwyg = "true";
defparam \mem[0][66] .power_up = "low";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][78] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_78_0),
	.prn(vcc));
defparam \mem[0][78] .is_wysiwyg = "true";
defparam \mem[0][78] .power_up = "low";

dffeas \mem[0][77] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_77_0),
	.prn(vcc));
defparam \mem[0][77] .is_wysiwyg = "true";
defparam \mem[0][77] .power_up = "low";

dffeas \mem[0][76] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_76_0),
	.prn(vcc));
defparam \mem[0][76] .is_wysiwyg = "true";
defparam \mem[0][76] .power_up = "low";

dffeas \mem[0][75] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_75_0),
	.prn(vcc));
defparam \mem[0][75] .is_wysiwyg = "true";
defparam \mem[0][75] .power_up = "low";

dffeas \mem[0][74] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_74_0),
	.prn(vcc));
defparam \mem[0][74] .is_wysiwyg = "true";
defparam \mem[0][74] .power_up = "low";

dffeas \mem[0][105] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_105_0),
	.prn(vcc));
defparam \mem[0][105] .is_wysiwyg = "true";
defparam \mem[0][105] .power_up = "low";

dffeas \mem[0][106] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_106_0),
	.prn(vcc));
defparam \mem[0][106] .is_wysiwyg = "true";
defparam \mem[0][106] .power_up = "low";

dffeas \mem[0][107] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_107_0),
	.prn(vcc));
defparam \mem[0][107] .is_wysiwyg = "true";
defparam \mem[0][107] .power_up = "low";

dffeas \mem[0][108] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_108_0),
	.prn(vcc));
defparam \mem[0][108] .is_wysiwyg = "true";
defparam \mem[0][108] .power_up = "low";

dffeas \mem[0][109] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_109_0),
	.prn(vcc));
defparam \mem[0][109] .is_wysiwyg = "true";
defparam \mem[0][109] .power_up = "low";

dffeas \mem[0][110] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_110_0),
	.prn(vcc));
defparam \mem[0][110] .is_wysiwyg = "true";
defparam \mem[0][110] .power_up = "low";

dffeas \mem[0][111] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_111_0),
	.prn(vcc));
defparam \mem[0][111] .is_wysiwyg = "true";
defparam \mem[0][111] .power_up = "low";

dffeas \mem[0][112] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_112_0),
	.prn(vcc));
defparam \mem[0][112] .is_wysiwyg = "true";
defparam \mem[0][112] .power_up = "low";

dffeas \mem[0][113] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_113_0),
	.prn(vcc));
defparam \mem[0][113] .is_wysiwyg = "true";
defparam \mem[0][113] .power_up = "low";

dffeas \mem[0][114] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_114_0),
	.prn(vcc));
defparam \mem[0][114] .is_wysiwyg = "true";
defparam \mem[0][114] .power_up = "low";

dffeas \mem[0][115] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_115_0),
	.prn(vcc));
defparam \mem[0][115] .is_wysiwyg = "true";
defparam \mem[0][115] .power_up = "low";

dffeas \mem[0][116] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_116_0),
	.prn(vcc));
defparam \mem[0][116] .is_wysiwyg = "true";
defparam \mem[0][116] .power_up = "low";

cyclonev_lcell_comb \write~0 (
	.dataa(!waitrequest_reset_override),
	.datab(!in_data_reg_69),
	.datac(!mem_used_1),
	.datad(!out_valid_reg),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'h0010001000100010;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \write~1 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!write),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write1),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~1 .extended_lut = "off";
defparam \write~1 .lut_mask = 64'h0202020202020202;
defparam \write~1 .shared_arith = "off";

cyclonev_lcell_comb \read~0 (
	.dataa(!h2f_RREADY_0),
	.datab(!empty),
	.datac(!last_packet_beat),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h4040404040404040;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!\read~0_combout ),
	.datad(!write1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'h5431543154315431;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][130] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][130]~q ),
	.prn(vcc));
defparam \mem[1][130] .is_wysiwyg = "true";
defparam \mem[1][130] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!mem_used_1),
	.datab(!nxt_out_eop),
	.datac(!\mem[1][130]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h2727272727272727;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!mem_used_0),
	.datab(!\read~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \always0~0 .shared_arith = "off";

dffeas \mem[1][69] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][69]~q ),
	.prn(vcc));
defparam \mem[1][69] .is_wysiwyg = "true";
defparam \mem[1][69] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!in_data_reg_69),
	.datab(!mem_used_1),
	.datac(!\mem[1][69]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h4747474747474747;
defparam \mem~1 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!\read~0_combout ),
	.datad(!write1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'h31FF31FF31FF31FF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem[1][78] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][78]~q ),
	.prn(vcc));
defparam \mem[1][78] .is_wysiwyg = "true";
defparam \mem[1][78] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_6),
	.datad(!\mem[1][78]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h0257025702570257;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[1][77] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][77]~q ),
	.prn(vcc));
defparam \mem[1][77] .is_wysiwyg = "true";
defparam \mem[1][77] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\mem[1][77]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h0257025702570257;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][76] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][76]~q ),
	.prn(vcc));
defparam \mem[1][76] .is_wysiwyg = "true";
defparam \mem[1][76] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!\mem[1][76]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h0257025702570257;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][75] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][75]~q ),
	.prn(vcc));
defparam \mem[1][75] .is_wysiwyg = "true";
defparam \mem[1][75] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\mem[1][75]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h0257025702570257;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][74] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][74]~q ),
	.prn(vcc));
defparam \mem[1][74] .is_wysiwyg = "true";
defparam \mem[1][74] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_byte_cnt_reg_2),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(!\mem[1][74]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h082A5D7F082A5D7F;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[1][105] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][105]~q ),
	.prn(vcc));
defparam \mem[1][105] .is_wysiwyg = "true";
defparam \mem[1][105] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][105]~q ),
	.datac(!in_data_reg_105),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[1][106] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][106]~q ),
	.prn(vcc));
defparam \mem[1][106] .is_wysiwyg = "true";
defparam \mem[1][106] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][106]~q ),
	.datac(!in_data_reg_106),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~8 .shared_arith = "off";

dffeas \mem[1][107] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][107]~q ),
	.prn(vcc));
defparam \mem[1][107] .is_wysiwyg = "true";
defparam \mem[1][107] .power_up = "low";

cyclonev_lcell_comb \mem~9 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][107]~q ),
	.datac(!in_data_reg_107),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~9 .extended_lut = "off";
defparam \mem~9 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~9 .shared_arith = "off";

dffeas \mem[1][108] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][108]~q ),
	.prn(vcc));
defparam \mem[1][108] .is_wysiwyg = "true";
defparam \mem[1][108] .power_up = "low";

cyclonev_lcell_comb \mem~10 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][108]~q ),
	.datac(!in_data_reg_108),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~10 .extended_lut = "off";
defparam \mem~10 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~10 .shared_arith = "off";

dffeas \mem[1][109] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][109]~q ),
	.prn(vcc));
defparam \mem[1][109] .is_wysiwyg = "true";
defparam \mem[1][109] .power_up = "low";

cyclonev_lcell_comb \mem~11 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][109]~q ),
	.datac(!in_data_reg_109),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~11 .extended_lut = "off";
defparam \mem~11 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~11 .shared_arith = "off";

dffeas \mem[1][110] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][110]~q ),
	.prn(vcc));
defparam \mem[1][110] .is_wysiwyg = "true";
defparam \mem[1][110] .power_up = "low";

cyclonev_lcell_comb \mem~12 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][110]~q ),
	.datac(!in_data_reg_110),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~12 .extended_lut = "off";
defparam \mem~12 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~12 .shared_arith = "off";

dffeas \mem[1][111] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][111]~q ),
	.prn(vcc));
defparam \mem[1][111] .is_wysiwyg = "true";
defparam \mem[1][111] .power_up = "low";

cyclonev_lcell_comb \mem~13 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][111]~q ),
	.datac(!in_data_reg_111),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~13 .extended_lut = "off";
defparam \mem~13 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~13 .shared_arith = "off";

dffeas \mem[1][112] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][112]~q ),
	.prn(vcc));
defparam \mem[1][112] .is_wysiwyg = "true";
defparam \mem[1][112] .power_up = "low";

cyclonev_lcell_comb \mem~14 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][112]~q ),
	.datac(!in_data_reg_112),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~14 .extended_lut = "off";
defparam \mem~14 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~14 .shared_arith = "off";

dffeas \mem[1][113] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][113]~q ),
	.prn(vcc));
defparam \mem[1][113] .is_wysiwyg = "true";
defparam \mem[1][113] .power_up = "low";

cyclonev_lcell_comb \mem~15 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][113]~q ),
	.datac(!in_data_reg_113),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~15 .extended_lut = "off";
defparam \mem~15 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~15 .shared_arith = "off";

dffeas \mem[1][114] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][114]~q ),
	.prn(vcc));
defparam \mem[1][114] .is_wysiwyg = "true";
defparam \mem[1][114] .power_up = "low";

cyclonev_lcell_comb \mem~16 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][114]~q ),
	.datac(!in_data_reg_114),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~16 .extended_lut = "off";
defparam \mem~16 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~16 .shared_arith = "off";

dffeas \mem[1][115] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][115]~q ),
	.prn(vcc));
defparam \mem[1][115] .is_wysiwyg = "true";
defparam \mem[1][115] .power_up = "low";

cyclonev_lcell_comb \mem~17 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][115]~q ),
	.datac(!in_data_reg_115),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~17 .extended_lut = "off";
defparam \mem~17 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~17 .shared_arith = "off";

dffeas \mem[1][116] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][116]~q ),
	.prn(vcc));
defparam \mem[1][116] .is_wysiwyg = "true";
defparam \mem[1][116] .power_up = "low";

cyclonev_lcell_comb \mem~18 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][116]~q ),
	.datac(!in_data_reg_116),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~18 .extended_lut = "off";
defparam \mem~18 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~18 .shared_arith = "off";

endmodule

module spw_babasu_altera_avalon_sc_fifo_4 (
	read_latency_shift_reg_0,
	mem_used_0,
	mem_129_0,
	mem_used_01,
	av_readdata_pre_0,
	always4,
	mem_0_0,
	av_readdata_pre_1,
	mem_1_0,
	av_readdata_pre_2,
	mem_2_0,
	av_readdata_pre_3,
	mem_3_0,
	av_readdata_pre_4,
	mem_4_0,
	av_readdata_pre_5,
	mem_5_0,
	av_readdata_pre_6,
	mem_6_0,
	av_readdata_pre_7,
	mem_7_0,
	av_readdata_pre_8,
	mem_8_0,
	reset,
	WideOr0,
	clk)/* synthesis synthesis_greybox=0 */;
input 	read_latency_shift_reg_0;
output 	mem_used_0;
input 	mem_129_0;
input 	mem_used_01;
input 	av_readdata_pre_0;
output 	always4;
output 	mem_0_0;
input 	av_readdata_pre_1;
output 	mem_1_0;
input 	av_readdata_pre_2;
output 	mem_2_0;
input 	av_readdata_pre_3;
output 	mem_3_0;
input 	av_readdata_pre_4;
output 	mem_4_0;
input 	av_readdata_pre_5;
output 	mem_5_0;
input 	av_readdata_pre_6;
output 	mem_6_0;
input 	av_readdata_pre_7;
output 	mem_7_0;
input 	av_readdata_pre_8;
output 	mem_8_0;
input 	reset;
input 	WideOr0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~q ;
wire \mem_used[0]~0_combout ;
wire \mem[1][0]~q ;
wire \mem~0_combout ;
wire \always0~0_combout ;
wire \mem[1][1]~q ;
wire \mem~1_combout ;
wire \mem[1][2]~q ;
wire \mem~2_combout ;
wire \mem[1][3]~q ;
wire \mem~3_combout ;
wire \mem[1][4]~q ;
wire \mem~4_combout ;
wire \mem[1][5]~q ;
wire \mem~5_combout ;
wire \mem[1][6]~q ;
wire \mem~6_combout ;
wire \mem[1][7]~q ;
wire \mem~7_combout ;
wire \mem[1][8]~q ;
wire \mem~8_combout ;


dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \always4~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always4),
	.sumout(),
	.cout(),
	.shareout());
defparam \always4~0 .extended_lut = "off";
defparam \always4~0 .lut_mask = 64'h4444444444444444;
defparam \always4~0 .shared_arith = "off";

dffeas \mem[0][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_0_0),
	.prn(vcc));
defparam \mem[0][0] .is_wysiwyg = "true";
defparam \mem[0][0] .power_up = "low";

dffeas \mem[0][1] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_1_0),
	.prn(vcc));
defparam \mem[0][1] .is_wysiwyg = "true";
defparam \mem[0][1] .power_up = "low";

dffeas \mem[0][2] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_2_0),
	.prn(vcc));
defparam \mem[0][2] .is_wysiwyg = "true";
defparam \mem[0][2] .power_up = "low";

dffeas \mem[0][3] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_3_0),
	.prn(vcc));
defparam \mem[0][3] .is_wysiwyg = "true";
defparam \mem[0][3] .power_up = "low";

dffeas \mem[0][4] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_4_0),
	.prn(vcc));
defparam \mem[0][4] .is_wysiwyg = "true";
defparam \mem[0][4] .power_up = "low";

dffeas \mem[0][5] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_5_0),
	.prn(vcc));
defparam \mem[0][5] .is_wysiwyg = "true";
defparam \mem[0][5] .power_up = "low";

dffeas \mem[0][6] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_6_0),
	.prn(vcc));
defparam \mem[0][6] .is_wysiwyg = "true";
defparam \mem[0][6] .power_up = "low";

dffeas \mem[0][7] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_7_0),
	.prn(vcc));
defparam \mem[0][7] .is_wysiwyg = "true";
defparam \mem[0][7] .power_up = "low";

dffeas \mem[0][8] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_8_0),
	.prn(vcc));
defparam \mem[0][8] .is_wysiwyg = "true";
defparam \mem[0][8] .power_up = "low";

cyclonev_lcell_comb \read~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_129_0),
	.datad(!mem_used_01),
	.datae(!WideOr0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h0000777000007770;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!\mem_used[1]~q ),
	.datad(!\read~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'h1F001F001F001F00;
defparam \mem_used[1]~1 .shared_arith = "off";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[1]~q ),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!\mem_used[1]~q ),
	.datad(!\read~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~0 .extended_lut = "off";
defparam \mem_used[0]~0 .lut_mask = 64'h731F731F731F731F;
defparam \mem_used[0]~0 .shared_arith = "off";

dffeas \mem[1][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][0]~q ),
	.prn(vcc));
defparam \mem[1][0] .is_wysiwyg = "true";
defparam \mem[1][0] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!av_readdata_pre_0),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h4747474747474747;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!mem_used_0),
	.datab(!\read~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \always0~0 .shared_arith = "off";

dffeas \mem[1][1] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][1]~q ),
	.prn(vcc));
defparam \mem[1][1] .is_wysiwyg = "true";
defparam \mem[1][1] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!av_readdata_pre_1),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h4747474747474747;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[1][2] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][2]~q ),
	.prn(vcc));
defparam \mem[1][2] .is_wysiwyg = "true";
defparam \mem[1][2] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!av_readdata_pre_2),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h4747474747474747;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[1][3] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][3]~q ),
	.prn(vcc));
defparam \mem[1][3] .is_wysiwyg = "true";
defparam \mem[1][3] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!av_readdata_pre_3),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h4747474747474747;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][4] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][4]~q ),
	.prn(vcc));
defparam \mem[1][4] .is_wysiwyg = "true";
defparam \mem[1][4] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!av_readdata_pre_4),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h4747474747474747;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][5] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][5]~q ),
	.prn(vcc));
defparam \mem[1][5] .is_wysiwyg = "true";
defparam \mem[1][5] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!av_readdata_pre_5),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][5]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h4747474747474747;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][6] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][6]~q ),
	.prn(vcc));
defparam \mem[1][6] .is_wysiwyg = "true";
defparam \mem[1][6] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!av_readdata_pre_6),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][6]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h4747474747474747;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[1][7] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][7]~q ),
	.prn(vcc));
defparam \mem[1][7] .is_wysiwyg = "true";
defparam \mem[1][7] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!av_readdata_pre_7),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h4747474747474747;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[1][8] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][8]~q ),
	.prn(vcc));
defparam \mem[1][8] .is_wysiwyg = "true";
defparam \mem[1][8] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!av_readdata_pre_8),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][8]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h4747474747474747;
defparam \mem~8 .shared_arith = "off";

endmodule

module spw_babasu_altera_avalon_sc_fifo_5 (
	out_valid_reg,
	mem_used_1,
	WideOr0,
	in_data_reg_68,
	stateST_UNCOMP_WR_SUBBURST,
	mem_129_0,
	mem_used_0,
	mem_68_0,
	mem_66_0,
	comb,
	mem_130_0,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	mem_105_0,
	mem_106_0,
	mem_107_0,
	mem_108_0,
	mem_109_0,
	mem_110_0,
	mem_111_0,
	mem_112_0,
	mem_113_0,
	mem_114_0,
	mem_115_0,
	mem_116_0,
	reset,
	nxt_out_eop,
	last_packet_beat,
	WideOr01,
	read,
	cp_ready,
	in_data_reg_69,
	rf_source_valid,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_6,
	sink_ready,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	clk)/* synthesis synthesis_greybox=0 */;
input 	out_valid_reg;
output 	mem_used_1;
input 	WideOr0;
input 	in_data_reg_68;
input 	stateST_UNCOMP_WR_SUBBURST;
output 	mem_129_0;
output 	mem_used_0;
output 	mem_68_0;
output 	mem_66_0;
input 	comb;
output 	mem_130_0;
output 	mem_78_0;
output 	mem_77_0;
output 	mem_76_0;
output 	mem_75_0;
output 	mem_74_0;
output 	mem_105_0;
output 	mem_106_0;
output 	mem_107_0;
output 	mem_108_0;
output 	mem_109_0;
output 	mem_110_0;
output 	mem_111_0;
output 	mem_112_0;
output 	mem_113_0;
output 	mem_114_0;
output 	mem_115_0;
output 	mem_116_0;
input 	reset;
input 	nxt_out_eop;
input 	last_packet_beat;
input 	WideOr01;
output 	read;
input 	cp_ready;
input 	in_data_reg_69;
input 	rf_source_valid;
input 	out_byte_cnt_reg_2;
input 	out_uncomp_byte_cnt_reg_3;
input 	out_uncomp_byte_cnt_reg_2;
input 	out_uncomp_byte_cnt_reg_4;
input 	out_uncomp_byte_cnt_reg_5;
input 	out_uncomp_byte_cnt_reg_6;
input 	sink_ready;
input 	in_data_reg_105;
input 	in_data_reg_106;
input 	in_data_reg_107;
input 	in_data_reg_108;
input 	in_data_reg_109;
input 	in_data_reg_110;
input 	in_data_reg_111;
input 	in_data_reg_112;
input 	in_data_reg_113;
input 	in_data_reg_114;
input 	in_data_reg_115;
input 	in_data_reg_116;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \write~0_combout ;
wire \mem_used[1]~0_combout ;
wire \mem[1][129]~q ;
wire \mem~20_combout ;
wire \always0~0_combout ;
wire \mem_used[0]~1_combout ;
wire \mem[1][68]~q ;
wire \mem~0_combout ;
wire \mem[1][69]~q ;
wire \mem~1_combout ;
wire \mem[1][130]~q ;
wire \mem~2_combout ;
wire \mem[1][78]~q ;
wire \mem~3_combout ;
wire \mem[1][77]~q ;
wire \mem~4_combout ;
wire \mem[1][76]~q ;
wire \mem~5_combout ;
wire \mem[1][75]~q ;
wire \mem~6_combout ;
wire \mem[1][74]~q ;
wire \mem~7_combout ;
wire \mem[1][105]~q ;
wire \mem~8_combout ;
wire \mem[1][106]~q ;
wire \mem~9_combout ;
wire \mem[1][107]~q ;
wire \mem~10_combout ;
wire \mem[1][108]~q ;
wire \mem~11_combout ;
wire \mem[1][109]~q ;
wire \mem~12_combout ;
wire \mem[1][110]~q ;
wire \mem~13_combout ;
wire \mem[1][111]~q ;
wire \mem~14_combout ;
wire \mem[1][112]~q ;
wire \mem~15_combout ;
wire \mem[1][113]~q ;
wire \mem~16_combout ;
wire \mem[1][114]~q ;
wire \mem~17_combout ;
wire \mem[1][115]~q ;
wire \mem~18_combout ;
wire \mem[1][116]~q ;
wire \mem~19_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][129] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_129_0),
	.prn(vcc));
defparam \mem[0][129] .is_wysiwyg = "true";
defparam \mem[0][129] .power_up = "low";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][68] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_68_0),
	.prn(vcc));
defparam \mem[0][68] .is_wysiwyg = "true";
defparam \mem[0][68] .power_up = "low";

dffeas \mem[0][66] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_66_0),
	.prn(vcc));
defparam \mem[0][66] .is_wysiwyg = "true";
defparam \mem[0][66] .power_up = "low";

dffeas \mem[0][130] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_130_0),
	.prn(vcc));
defparam \mem[0][130] .is_wysiwyg = "true";
defparam \mem[0][130] .power_up = "low";

dffeas \mem[0][78] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_78_0),
	.prn(vcc));
defparam \mem[0][78] .is_wysiwyg = "true";
defparam \mem[0][78] .power_up = "low";

dffeas \mem[0][77] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_77_0),
	.prn(vcc));
defparam \mem[0][77] .is_wysiwyg = "true";
defparam \mem[0][77] .power_up = "low";

dffeas \mem[0][76] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_76_0),
	.prn(vcc));
defparam \mem[0][76] .is_wysiwyg = "true";
defparam \mem[0][76] .power_up = "low";

dffeas \mem[0][75] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_75_0),
	.prn(vcc));
defparam \mem[0][75] .is_wysiwyg = "true";
defparam \mem[0][75] .power_up = "low";

dffeas \mem[0][74] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_74_0),
	.prn(vcc));
defparam \mem[0][74] .is_wysiwyg = "true";
defparam \mem[0][74] .power_up = "low";

dffeas \mem[0][105] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_105_0),
	.prn(vcc));
defparam \mem[0][105] .is_wysiwyg = "true";
defparam \mem[0][105] .power_up = "low";

dffeas \mem[0][106] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_106_0),
	.prn(vcc));
defparam \mem[0][106] .is_wysiwyg = "true";
defparam \mem[0][106] .power_up = "low";

dffeas \mem[0][107] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_107_0),
	.prn(vcc));
defparam \mem[0][107] .is_wysiwyg = "true";
defparam \mem[0][107] .power_up = "low";

dffeas \mem[0][108] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_108_0),
	.prn(vcc));
defparam \mem[0][108] .is_wysiwyg = "true";
defparam \mem[0][108] .power_up = "low";

dffeas \mem[0][109] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_109_0),
	.prn(vcc));
defparam \mem[0][109] .is_wysiwyg = "true";
defparam \mem[0][109] .power_up = "low";

dffeas \mem[0][110] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_110_0),
	.prn(vcc));
defparam \mem[0][110] .is_wysiwyg = "true";
defparam \mem[0][110] .power_up = "low";

dffeas \mem[0][111] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_111_0),
	.prn(vcc));
defparam \mem[0][111] .is_wysiwyg = "true";
defparam \mem[0][111] .power_up = "low";

dffeas \mem[0][112] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_112_0),
	.prn(vcc));
defparam \mem[0][112] .is_wysiwyg = "true";
defparam \mem[0][112] .power_up = "low";

dffeas \mem[0][113] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_113_0),
	.prn(vcc));
defparam \mem[0][113] .is_wysiwyg = "true";
defparam \mem[0][113] .power_up = "low";

dffeas \mem[0][114] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_114_0),
	.prn(vcc));
defparam \mem[0][114] .is_wysiwyg = "true";
defparam \mem[0][114] .power_up = "low";

dffeas \mem[0][115] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_115_0),
	.prn(vcc));
defparam \mem[0][115] .is_wysiwyg = "true";
defparam \mem[0][115] .power_up = "low";

dffeas \mem[0][116] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_116_0),
	.prn(vcc));
defparam \mem[0][116] .is_wysiwyg = "true";
defparam \mem[0][116] .power_up = "low";

cyclonev_lcell_comb \read~0 (
	.dataa(!comb),
	.datab(!WideOr01),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h1111111111111111;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \write~0 (
	.dataa(!mem_used_1),
	.datab(!WideOr0),
	.datac(!cp_ready),
	.datad(!rf_source_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'h008A008A008A008A;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!last_packet_beat),
	.datad(!read),
	.datae(!\write~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'h5505335355053353;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][129] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][129]~q ),
	.prn(vcc));
defparam \mem[1][129] .is_wysiwyg = "true";
defparam \mem[1][129] .power_up = "low";

cyclonev_lcell_comb \mem~20 (
	.dataa(!WideOr0),
	.datab(!out_valid_reg),
	.datac(!\mem[1][129]~q ),
	.datad(!in_data_reg_68),
	.datae(!mem_used_1),
	.dataf(!nxt_out_eop),
	.datag(!in_data_reg_69),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~20 .extended_lut = "on";
defparam \mem~20 .lut_mask = 64'h02020F0F02330F0F;
defparam \mem~20 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!mem_used_0),
	.datab(!sink_ready),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!\write~0_combout ),
	.datad(!sink_ready),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'h3F1F3F1F3F1F3F1F;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem[1][68] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][68]~q ),
	.prn(vcc));
defparam \mem[1][68] .is_wysiwyg = "true";
defparam \mem[1][68] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!mem_used_1),
	.datab(!in_data_reg_68),
	.datac(!\mem[1][68]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h2727272727272727;
defparam \mem~0 .shared_arith = "off";

dffeas \mem[1][69] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][69]~q ),
	.prn(vcc));
defparam \mem[1][69] .is_wysiwyg = "true";
defparam \mem[1][69] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!mem_used_1),
	.datab(!in_data_reg_69),
	.datac(!\mem[1][69]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h2727272727272727;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[1][130] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][130]~q ),
	.prn(vcc));
defparam \mem[1][130] .is_wysiwyg = "true";
defparam \mem[1][130] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!mem_used_1),
	.datab(!nxt_out_eop),
	.datac(!\mem[1][130]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h2727272727272727;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[1][78] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][78]~q ),
	.prn(vcc));
defparam \mem[1][78] .is_wysiwyg = "true";
defparam \mem[1][78] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_6),
	.datad(!\mem[1][78]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h0257025702570257;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][77] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][77]~q ),
	.prn(vcc));
defparam \mem[1][77] .is_wysiwyg = "true";
defparam \mem[1][77] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\mem[1][77]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h0257025702570257;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][76] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][76]~q ),
	.prn(vcc));
defparam \mem[1][76] .is_wysiwyg = "true";
defparam \mem[1][76] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!\mem[1][76]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h0257025702570257;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][75] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][75]~q ),
	.prn(vcc));
defparam \mem[1][75] .is_wysiwyg = "true";
defparam \mem[1][75] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\mem[1][75]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h0257025702570257;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[1][74] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][74]~q ),
	.prn(vcc));
defparam \mem[1][74] .is_wysiwyg = "true";
defparam \mem[1][74] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_byte_cnt_reg_2),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(!\mem[1][74]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h082A5D7F082A5D7F;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[1][105] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][105]~q ),
	.prn(vcc));
defparam \mem[1][105] .is_wysiwyg = "true";
defparam \mem[1][105] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][105]~q ),
	.datac(!in_data_reg_105),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~8 .shared_arith = "off";

dffeas \mem[1][106] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][106]~q ),
	.prn(vcc));
defparam \mem[1][106] .is_wysiwyg = "true";
defparam \mem[1][106] .power_up = "low";

cyclonev_lcell_comb \mem~9 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][106]~q ),
	.datac(!in_data_reg_106),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~9 .extended_lut = "off";
defparam \mem~9 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~9 .shared_arith = "off";

dffeas \mem[1][107] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][107]~q ),
	.prn(vcc));
defparam \mem[1][107] .is_wysiwyg = "true";
defparam \mem[1][107] .power_up = "low";

cyclonev_lcell_comb \mem~10 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][107]~q ),
	.datac(!in_data_reg_107),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~10 .extended_lut = "off";
defparam \mem~10 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~10 .shared_arith = "off";

dffeas \mem[1][108] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][108]~q ),
	.prn(vcc));
defparam \mem[1][108] .is_wysiwyg = "true";
defparam \mem[1][108] .power_up = "low";

cyclonev_lcell_comb \mem~11 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][108]~q ),
	.datac(!in_data_reg_108),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~11 .extended_lut = "off";
defparam \mem~11 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~11 .shared_arith = "off";

dffeas \mem[1][109] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][109]~q ),
	.prn(vcc));
defparam \mem[1][109] .is_wysiwyg = "true";
defparam \mem[1][109] .power_up = "low";

cyclonev_lcell_comb \mem~12 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][109]~q ),
	.datac(!in_data_reg_109),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~12 .extended_lut = "off";
defparam \mem~12 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~12 .shared_arith = "off";

dffeas \mem[1][110] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][110]~q ),
	.prn(vcc));
defparam \mem[1][110] .is_wysiwyg = "true";
defparam \mem[1][110] .power_up = "low";

cyclonev_lcell_comb \mem~13 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][110]~q ),
	.datac(!in_data_reg_110),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~13 .extended_lut = "off";
defparam \mem~13 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~13 .shared_arith = "off";

dffeas \mem[1][111] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][111]~q ),
	.prn(vcc));
defparam \mem[1][111] .is_wysiwyg = "true";
defparam \mem[1][111] .power_up = "low";

cyclonev_lcell_comb \mem~14 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][111]~q ),
	.datac(!in_data_reg_111),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~14 .extended_lut = "off";
defparam \mem~14 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~14 .shared_arith = "off";

dffeas \mem[1][112] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][112]~q ),
	.prn(vcc));
defparam \mem[1][112] .is_wysiwyg = "true";
defparam \mem[1][112] .power_up = "low";

cyclonev_lcell_comb \mem~15 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][112]~q ),
	.datac(!in_data_reg_112),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~15 .extended_lut = "off";
defparam \mem~15 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~15 .shared_arith = "off";

dffeas \mem[1][113] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][113]~q ),
	.prn(vcc));
defparam \mem[1][113] .is_wysiwyg = "true";
defparam \mem[1][113] .power_up = "low";

cyclonev_lcell_comb \mem~16 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][113]~q ),
	.datac(!in_data_reg_113),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~16 .extended_lut = "off";
defparam \mem~16 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~16 .shared_arith = "off";

dffeas \mem[1][114] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][114]~q ),
	.prn(vcc));
defparam \mem[1][114] .is_wysiwyg = "true";
defparam \mem[1][114] .power_up = "low";

cyclonev_lcell_comb \mem~17 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][114]~q ),
	.datac(!in_data_reg_114),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~17 .extended_lut = "off";
defparam \mem~17 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~17 .shared_arith = "off";

dffeas \mem[1][115] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][115]~q ),
	.prn(vcc));
defparam \mem[1][115] .is_wysiwyg = "true";
defparam \mem[1][115] .power_up = "low";

cyclonev_lcell_comb \mem~18 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][115]~q ),
	.datac(!in_data_reg_115),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~18 .extended_lut = "off";
defparam \mem~18 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~18 .shared_arith = "off";

dffeas \mem[1][116] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][116]~q ),
	.prn(vcc));
defparam \mem[1][116] .is_wysiwyg = "true";
defparam \mem[1][116] .power_up = "low";

cyclonev_lcell_comb \mem~19 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][116]~q ),
	.datac(!in_data_reg_116),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~19 .extended_lut = "off";
defparam \mem~19 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~19 .shared_arith = "off";

endmodule

module spw_babasu_altera_avalon_sc_fifo_6 (
	h2f_RREADY_0,
	read_latency_shift_reg_0,
	mem_used_0,
	empty1,
	av_readdata_pre_0,
	mem_0_0,
	mem_1_0,
	av_readdata_pre_1,
	mem_2_0,
	av_readdata_pre_2,
	mem_3_0,
	av_readdata_pre_3,
	mem_4_0,
	av_readdata_pre_4,
	mem_5_0,
	av_readdata_pre_5,
	mem_6_0,
	av_readdata_pre_6,
	mem_7_0,
	av_readdata_pre_7,
	mem_8_0,
	av_readdata_pre_8,
	reset,
	clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_RREADY_0;
input 	read_latency_shift_reg_0;
output 	mem_used_0;
output 	empty1;
input 	av_readdata_pre_0;
output 	mem_0_0;
output 	mem_1_0;
input 	av_readdata_pre_1;
output 	mem_2_0;
input 	av_readdata_pre_2;
output 	mem_3_0;
input 	av_readdata_pre_3;
output 	mem_4_0;
input 	av_readdata_pre_4;
output 	mem_5_0;
input 	av_readdata_pre_5;
output 	mem_6_0;
input 	av_readdata_pre_6;
output 	mem_7_0;
input 	av_readdata_pre_7;
output 	mem_8_0;
input 	av_readdata_pre_8;
input 	reset;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[1]~1_combout ;
wire \mem_used[1]~q ;
wire \mem_used[0]~0_combout ;
wire \mem[1][0]~q ;
wire \mem~0_combout ;
wire \always0~0_combout ;
wire \mem[1][1]~q ;
wire \mem~1_combout ;
wire \mem[1][2]~q ;
wire \mem~2_combout ;
wire \mem[1][3]~q ;
wire \mem~3_combout ;
wire \mem[1][4]~q ;
wire \mem~4_combout ;
wire \mem[1][5]~q ;
wire \mem~5_combout ;
wire \mem[1][6]~q ;
wire \mem~6_combout ;
wire \mem[1][7]~q ;
wire \mem~7_combout ;
wire \mem[1][8]~q ;
wire \mem~8_combout ;


dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb empty(
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(empty1),
	.sumout(),
	.cout(),
	.shareout());
defparam empty.extended_lut = "off";
defparam empty.lut_mask = 64'h8888888888888888;
defparam empty.shared_arith = "off";

dffeas \mem[0][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_0_0),
	.prn(vcc));
defparam \mem[0][0] .is_wysiwyg = "true";
defparam \mem[0][0] .power_up = "low";

dffeas \mem[0][1] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_1_0),
	.prn(vcc));
defparam \mem[0][1] .is_wysiwyg = "true";
defparam \mem[0][1] .power_up = "low";

dffeas \mem[0][2] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_2_0),
	.prn(vcc));
defparam \mem[0][2] .is_wysiwyg = "true";
defparam \mem[0][2] .power_up = "low";

dffeas \mem[0][3] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_3_0),
	.prn(vcc));
defparam \mem[0][3] .is_wysiwyg = "true";
defparam \mem[0][3] .power_up = "low";

dffeas \mem[0][4] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_4_0),
	.prn(vcc));
defparam \mem[0][4] .is_wysiwyg = "true";
defparam \mem[0][4] .power_up = "low";

dffeas \mem[0][5] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_5_0),
	.prn(vcc));
defparam \mem[0][5] .is_wysiwyg = "true";
defparam \mem[0][5] .power_up = "low";

dffeas \mem[0][6] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_6_0),
	.prn(vcc));
defparam \mem[0][6] .is_wysiwyg = "true";
defparam \mem[0][6] .power_up = "low";

dffeas \mem[0][7] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_7_0),
	.prn(vcc));
defparam \mem[0][7] .is_wysiwyg = "true";
defparam \mem[0][7] .power_up = "low";

dffeas \mem[0][8] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_8_0),
	.prn(vcc));
defparam \mem[0][8] .is_wysiwyg = "true";
defparam \mem[0][8] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!h2f_RREADY_0),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem_used[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'h02EA02EA02EA02EA;
defparam \mem_used[1]~1 .shared_arith = "off";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[1]~q ),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~0 (
	.dataa(!h2f_RREADY_0),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem_used[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~0 .extended_lut = "off";
defparam \mem_used[0]~0 .lut_mask = 64'h2B1F2B1F2B1F2B1F;
defparam \mem_used[0]~0 .shared_arith = "off";

dffeas \mem[1][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][0]~q ),
	.prn(vcc));
defparam \mem[1][0] .is_wysiwyg = "true";
defparam \mem[1][0] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!av_readdata_pre_0),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h4747474747474747;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!h2f_RREADY_0),
	.datab(!mem_used_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \always0~0 .shared_arith = "off";

dffeas \mem[1][1] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][1]~q ),
	.prn(vcc));
defparam \mem[1][1] .is_wysiwyg = "true";
defparam \mem[1][1] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!av_readdata_pre_1),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h4747474747474747;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[1][2] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][2]~q ),
	.prn(vcc));
defparam \mem[1][2] .is_wysiwyg = "true";
defparam \mem[1][2] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!av_readdata_pre_2),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h4747474747474747;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[1][3] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][3]~q ),
	.prn(vcc));
defparam \mem[1][3] .is_wysiwyg = "true";
defparam \mem[1][3] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!av_readdata_pre_3),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h4747474747474747;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][4] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][4]~q ),
	.prn(vcc));
defparam \mem[1][4] .is_wysiwyg = "true";
defparam \mem[1][4] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!av_readdata_pre_4),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h4747474747474747;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][5] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][5]~q ),
	.prn(vcc));
defparam \mem[1][5] .is_wysiwyg = "true";
defparam \mem[1][5] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!av_readdata_pre_5),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][5]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h4747474747474747;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][6] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][6]~q ),
	.prn(vcc));
defparam \mem[1][6] .is_wysiwyg = "true";
defparam \mem[1][6] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!av_readdata_pre_6),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][6]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h4747474747474747;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[1][7] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][7]~q ),
	.prn(vcc));
defparam \mem[1][7] .is_wysiwyg = "true";
defparam \mem[1][7] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!av_readdata_pre_7),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h4747474747474747;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[1][8] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][8]~q ),
	.prn(vcc));
defparam \mem[1][8] .is_wysiwyg = "true";
defparam \mem[1][8] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!av_readdata_pre_8),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][8]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h4747474747474747;
defparam \mem~8 .shared_arith = "off";

endmodule

module spw_babasu_altera_avalon_sc_fifo_7 (
	h2f_RREADY_0,
	mem_used_1,
	waitrequest_reset_override,
	in_data_reg_69,
	wait_latency_counter_1,
	wait_latency_counter_0,
	nxt_out_eop,
	out_valid_reg,
	stateST_UNCOMP_WR_SUBBURST,
	mem_130_0,
	empty,
	mem_66_0,
	mem_used_0,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	mem_105_0,
	mem_106_0,
	mem_107_0,
	mem_108_0,
	mem_109_0,
	mem_110_0,
	mem_111_0,
	mem_112_0,
	mem_113_0,
	mem_114_0,
	mem_115_0,
	mem_116_0,
	reset,
	last_packet_beat,
	write,
	write1,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_6,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_RREADY_0;
output 	mem_used_1;
input 	waitrequest_reset_override;
input 	in_data_reg_69;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	nxt_out_eop;
input 	out_valid_reg;
input 	stateST_UNCOMP_WR_SUBBURST;
output 	mem_130_0;
input 	empty;
output 	mem_66_0;
output 	mem_used_0;
output 	mem_78_0;
output 	mem_77_0;
output 	mem_76_0;
output 	mem_75_0;
output 	mem_74_0;
output 	mem_105_0;
output 	mem_106_0;
output 	mem_107_0;
output 	mem_108_0;
output 	mem_109_0;
output 	mem_110_0;
output 	mem_111_0;
output 	mem_112_0;
output 	mem_113_0;
output 	mem_114_0;
output 	mem_115_0;
output 	mem_116_0;
input 	reset;
input 	last_packet_beat;
output 	write;
output 	write1;
input 	out_byte_cnt_reg_2;
input 	out_uncomp_byte_cnt_reg_6;
input 	out_uncomp_byte_cnt_reg_5;
input 	out_uncomp_byte_cnt_reg_4;
input 	out_uncomp_byte_cnt_reg_3;
input 	out_uncomp_byte_cnt_reg_2;
input 	in_data_reg_105;
input 	in_data_reg_106;
input 	in_data_reg_107;
input 	in_data_reg_108;
input 	in_data_reg_109;
input 	in_data_reg_110;
input 	in_data_reg_111;
input 	in_data_reg_112;
input 	in_data_reg_113;
input 	in_data_reg_114;
input 	in_data_reg_115;
input 	in_data_reg_116;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read~0_combout ;
wire \mem_used[1]~0_combout ;
wire \mem[1][130]~q ;
wire \mem~0_combout ;
wire \always0~0_combout ;
wire \mem[1][69]~q ;
wire \mem~1_combout ;
wire \mem_used[0]~1_combout ;
wire \mem[1][78]~q ;
wire \mem~2_combout ;
wire \mem[1][77]~q ;
wire \mem~3_combout ;
wire \mem[1][76]~q ;
wire \mem~4_combout ;
wire \mem[1][75]~q ;
wire \mem~5_combout ;
wire \mem[1][74]~q ;
wire \mem~6_combout ;
wire \mem[1][105]~q ;
wire \mem~7_combout ;
wire \mem[1][106]~q ;
wire \mem~8_combout ;
wire \mem[1][107]~q ;
wire \mem~9_combout ;
wire \mem[1][108]~q ;
wire \mem~10_combout ;
wire \mem[1][109]~q ;
wire \mem~11_combout ;
wire \mem[1][110]~q ;
wire \mem~12_combout ;
wire \mem[1][111]~q ;
wire \mem~13_combout ;
wire \mem[1][112]~q ;
wire \mem~14_combout ;
wire \mem[1][113]~q ;
wire \mem~15_combout ;
wire \mem[1][114]~q ;
wire \mem~16_combout ;
wire \mem[1][115]~q ;
wire \mem~17_combout ;
wire \mem[1][116]~q ;
wire \mem~18_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][130] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_130_0),
	.prn(vcc));
defparam \mem[0][130] .is_wysiwyg = "true";
defparam \mem[0][130] .power_up = "low";

dffeas \mem[0][66] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_66_0),
	.prn(vcc));
defparam \mem[0][66] .is_wysiwyg = "true";
defparam \mem[0][66] .power_up = "low";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][78] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_78_0),
	.prn(vcc));
defparam \mem[0][78] .is_wysiwyg = "true";
defparam \mem[0][78] .power_up = "low";

dffeas \mem[0][77] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_77_0),
	.prn(vcc));
defparam \mem[0][77] .is_wysiwyg = "true";
defparam \mem[0][77] .power_up = "low";

dffeas \mem[0][76] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_76_0),
	.prn(vcc));
defparam \mem[0][76] .is_wysiwyg = "true";
defparam \mem[0][76] .power_up = "low";

dffeas \mem[0][75] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_75_0),
	.prn(vcc));
defparam \mem[0][75] .is_wysiwyg = "true";
defparam \mem[0][75] .power_up = "low";

dffeas \mem[0][74] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_74_0),
	.prn(vcc));
defparam \mem[0][74] .is_wysiwyg = "true";
defparam \mem[0][74] .power_up = "low";

dffeas \mem[0][105] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_105_0),
	.prn(vcc));
defparam \mem[0][105] .is_wysiwyg = "true";
defparam \mem[0][105] .power_up = "low";

dffeas \mem[0][106] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_106_0),
	.prn(vcc));
defparam \mem[0][106] .is_wysiwyg = "true";
defparam \mem[0][106] .power_up = "low";

dffeas \mem[0][107] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_107_0),
	.prn(vcc));
defparam \mem[0][107] .is_wysiwyg = "true";
defparam \mem[0][107] .power_up = "low";

dffeas \mem[0][108] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_108_0),
	.prn(vcc));
defparam \mem[0][108] .is_wysiwyg = "true";
defparam \mem[0][108] .power_up = "low";

dffeas \mem[0][109] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_109_0),
	.prn(vcc));
defparam \mem[0][109] .is_wysiwyg = "true";
defparam \mem[0][109] .power_up = "low";

dffeas \mem[0][110] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_110_0),
	.prn(vcc));
defparam \mem[0][110] .is_wysiwyg = "true";
defparam \mem[0][110] .power_up = "low";

dffeas \mem[0][111] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_111_0),
	.prn(vcc));
defparam \mem[0][111] .is_wysiwyg = "true";
defparam \mem[0][111] .power_up = "low";

dffeas \mem[0][112] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_112_0),
	.prn(vcc));
defparam \mem[0][112] .is_wysiwyg = "true";
defparam \mem[0][112] .power_up = "low";

dffeas \mem[0][113] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_113_0),
	.prn(vcc));
defparam \mem[0][113] .is_wysiwyg = "true";
defparam \mem[0][113] .power_up = "low";

dffeas \mem[0][114] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_114_0),
	.prn(vcc));
defparam \mem[0][114] .is_wysiwyg = "true";
defparam \mem[0][114] .power_up = "low";

dffeas \mem[0][115] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_115_0),
	.prn(vcc));
defparam \mem[0][115] .is_wysiwyg = "true";
defparam \mem[0][115] .power_up = "low";

dffeas \mem[0][116] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_116_0),
	.prn(vcc));
defparam \mem[0][116] .is_wysiwyg = "true";
defparam \mem[0][116] .power_up = "low";

cyclonev_lcell_comb \write~0 (
	.dataa(!waitrequest_reset_override),
	.datab(!in_data_reg_69),
	.datac(!mem_used_1),
	.datad(!out_valid_reg),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'h0010001000100010;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \write~1 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!write),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write1),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~1 .extended_lut = "off";
defparam \write~1 .lut_mask = 64'h0202020202020202;
defparam \write~1 .shared_arith = "off";

cyclonev_lcell_comb \read~0 (
	.dataa(!h2f_RREADY_0),
	.datab(!empty),
	.datac(!last_packet_beat),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h4040404040404040;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!\read~0_combout ),
	.datad(!write1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'h5431543154315431;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][130] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][130]~q ),
	.prn(vcc));
defparam \mem[1][130] .is_wysiwyg = "true";
defparam \mem[1][130] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!mem_used_1),
	.datab(!nxt_out_eop),
	.datac(!\mem[1][130]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h2727272727272727;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!mem_used_0),
	.datab(!\read~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \always0~0 .shared_arith = "off";

dffeas \mem[1][69] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][69]~q ),
	.prn(vcc));
defparam \mem[1][69] .is_wysiwyg = "true";
defparam \mem[1][69] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!in_data_reg_69),
	.datab(!mem_used_1),
	.datac(!\mem[1][69]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h4747474747474747;
defparam \mem~1 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!\read~0_combout ),
	.datad(!write1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'h31FF31FF31FF31FF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem[1][78] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][78]~q ),
	.prn(vcc));
defparam \mem[1][78] .is_wysiwyg = "true";
defparam \mem[1][78] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_6),
	.datad(!\mem[1][78]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h0257025702570257;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[1][77] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][77]~q ),
	.prn(vcc));
defparam \mem[1][77] .is_wysiwyg = "true";
defparam \mem[1][77] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\mem[1][77]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h0257025702570257;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][76] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][76]~q ),
	.prn(vcc));
defparam \mem[1][76] .is_wysiwyg = "true";
defparam \mem[1][76] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!\mem[1][76]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h0257025702570257;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][75] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][75]~q ),
	.prn(vcc));
defparam \mem[1][75] .is_wysiwyg = "true";
defparam \mem[1][75] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\mem[1][75]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h0257025702570257;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][74] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][74]~q ),
	.prn(vcc));
defparam \mem[1][74] .is_wysiwyg = "true";
defparam \mem[1][74] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_byte_cnt_reg_2),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(!\mem[1][74]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h082A5D7F082A5D7F;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[1][105] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][105]~q ),
	.prn(vcc));
defparam \mem[1][105] .is_wysiwyg = "true";
defparam \mem[1][105] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][105]~q ),
	.datac(!in_data_reg_105),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[1][106] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][106]~q ),
	.prn(vcc));
defparam \mem[1][106] .is_wysiwyg = "true";
defparam \mem[1][106] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][106]~q ),
	.datac(!in_data_reg_106),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~8 .shared_arith = "off";

dffeas \mem[1][107] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][107]~q ),
	.prn(vcc));
defparam \mem[1][107] .is_wysiwyg = "true";
defparam \mem[1][107] .power_up = "low";

cyclonev_lcell_comb \mem~9 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][107]~q ),
	.datac(!in_data_reg_107),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~9 .extended_lut = "off";
defparam \mem~9 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~9 .shared_arith = "off";

dffeas \mem[1][108] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][108]~q ),
	.prn(vcc));
defparam \mem[1][108] .is_wysiwyg = "true";
defparam \mem[1][108] .power_up = "low";

cyclonev_lcell_comb \mem~10 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][108]~q ),
	.datac(!in_data_reg_108),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~10 .extended_lut = "off";
defparam \mem~10 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~10 .shared_arith = "off";

dffeas \mem[1][109] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][109]~q ),
	.prn(vcc));
defparam \mem[1][109] .is_wysiwyg = "true";
defparam \mem[1][109] .power_up = "low";

cyclonev_lcell_comb \mem~11 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][109]~q ),
	.datac(!in_data_reg_109),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~11 .extended_lut = "off";
defparam \mem~11 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~11 .shared_arith = "off";

dffeas \mem[1][110] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][110]~q ),
	.prn(vcc));
defparam \mem[1][110] .is_wysiwyg = "true";
defparam \mem[1][110] .power_up = "low";

cyclonev_lcell_comb \mem~12 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][110]~q ),
	.datac(!in_data_reg_110),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~12 .extended_lut = "off";
defparam \mem~12 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~12 .shared_arith = "off";

dffeas \mem[1][111] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][111]~q ),
	.prn(vcc));
defparam \mem[1][111] .is_wysiwyg = "true";
defparam \mem[1][111] .power_up = "low";

cyclonev_lcell_comb \mem~13 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][111]~q ),
	.datac(!in_data_reg_111),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~13 .extended_lut = "off";
defparam \mem~13 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~13 .shared_arith = "off";

dffeas \mem[1][112] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][112]~q ),
	.prn(vcc));
defparam \mem[1][112] .is_wysiwyg = "true";
defparam \mem[1][112] .power_up = "low";

cyclonev_lcell_comb \mem~14 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][112]~q ),
	.datac(!in_data_reg_112),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~14 .extended_lut = "off";
defparam \mem~14 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~14 .shared_arith = "off";

dffeas \mem[1][113] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][113]~q ),
	.prn(vcc));
defparam \mem[1][113] .is_wysiwyg = "true";
defparam \mem[1][113] .power_up = "low";

cyclonev_lcell_comb \mem~15 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][113]~q ),
	.datac(!in_data_reg_113),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~15 .extended_lut = "off";
defparam \mem~15 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~15 .shared_arith = "off";

dffeas \mem[1][114] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][114]~q ),
	.prn(vcc));
defparam \mem[1][114] .is_wysiwyg = "true";
defparam \mem[1][114] .power_up = "low";

cyclonev_lcell_comb \mem~16 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][114]~q ),
	.datac(!in_data_reg_114),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~16 .extended_lut = "off";
defparam \mem~16 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~16 .shared_arith = "off";

dffeas \mem[1][115] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][115]~q ),
	.prn(vcc));
defparam \mem[1][115] .is_wysiwyg = "true";
defparam \mem[1][115] .power_up = "low";

cyclonev_lcell_comb \mem~17 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][115]~q ),
	.datac(!in_data_reg_115),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~17 .extended_lut = "off";
defparam \mem~17 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~17 .shared_arith = "off";

dffeas \mem[1][116] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][116]~q ),
	.prn(vcc));
defparam \mem[1][116] .is_wysiwyg = "true";
defparam \mem[1][116] .power_up = "low";

cyclonev_lcell_comb \mem~18 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][116]~q ),
	.datac(!in_data_reg_116),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~18 .extended_lut = "off";
defparam \mem~18 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~18 .shared_arith = "off";

endmodule

module spw_babasu_altera_avalon_sc_fifo_8 (
	h2f_RREADY_0,
	read_latency_shift_reg_0,
	mem_used_0,
	empty1,
	av_readdata_pre_0,
	mem_0_0,
	mem_1_0,
	av_readdata_pre_1,
	mem_2_0,
	av_readdata_pre_2,
	av_readdata_pre_3,
	mem_3_0,
	av_readdata_pre_4,
	mem_4_0,
	av_readdata_pre_5,
	mem_5_0,
	av_readdata_pre_6,
	mem_6_0,
	av_readdata_pre_7,
	mem_7_0,
	mem_8_0,
	av_readdata_pre_8,
	mem_9_0,
	av_readdata_pre_9,
	mem_10_0,
	av_readdata_pre_10,
	reset,
	clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_RREADY_0;
input 	read_latency_shift_reg_0;
output 	mem_used_0;
output 	empty1;
input 	av_readdata_pre_0;
output 	mem_0_0;
output 	mem_1_0;
input 	av_readdata_pre_1;
output 	mem_2_0;
input 	av_readdata_pre_2;
input 	av_readdata_pre_3;
output 	mem_3_0;
input 	av_readdata_pre_4;
output 	mem_4_0;
input 	av_readdata_pre_5;
output 	mem_5_0;
input 	av_readdata_pre_6;
output 	mem_6_0;
input 	av_readdata_pre_7;
output 	mem_7_0;
output 	mem_8_0;
input 	av_readdata_pre_8;
output 	mem_9_0;
input 	av_readdata_pre_9;
output 	mem_10_0;
input 	av_readdata_pre_10;
input 	reset;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[1]~1_combout ;
wire \mem_used[1]~q ;
wire \mem_used[0]~0_combout ;
wire \mem[1][0]~q ;
wire \mem~0_combout ;
wire \always0~0_combout ;
wire \mem[1][1]~q ;
wire \mem~1_combout ;
wire \mem[1][2]~q ;
wire \mem~2_combout ;
wire \mem[1][3]~q ;
wire \mem~3_combout ;
wire \mem[1][4]~q ;
wire \mem~4_combout ;
wire \mem[1][5]~q ;
wire \mem~5_combout ;
wire \mem[1][6]~q ;
wire \mem~6_combout ;
wire \mem[1][7]~q ;
wire \mem~7_combout ;
wire \mem[1][8]~q ;
wire \mem~8_combout ;
wire \mem[1][9]~q ;
wire \mem~9_combout ;
wire \mem[1][10]~q ;
wire \mem~10_combout ;


dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb empty(
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(empty1),
	.sumout(),
	.cout(),
	.shareout());
defparam empty.extended_lut = "off";
defparam empty.lut_mask = 64'h8888888888888888;
defparam empty.shared_arith = "off";

dffeas \mem[0][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_0_0),
	.prn(vcc));
defparam \mem[0][0] .is_wysiwyg = "true";
defparam \mem[0][0] .power_up = "low";

dffeas \mem[0][1] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_1_0),
	.prn(vcc));
defparam \mem[0][1] .is_wysiwyg = "true";
defparam \mem[0][1] .power_up = "low";

dffeas \mem[0][2] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_2_0),
	.prn(vcc));
defparam \mem[0][2] .is_wysiwyg = "true";
defparam \mem[0][2] .power_up = "low";

dffeas \mem[0][3] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_3_0),
	.prn(vcc));
defparam \mem[0][3] .is_wysiwyg = "true";
defparam \mem[0][3] .power_up = "low";

dffeas \mem[0][4] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_4_0),
	.prn(vcc));
defparam \mem[0][4] .is_wysiwyg = "true";
defparam \mem[0][4] .power_up = "low";

dffeas \mem[0][5] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_5_0),
	.prn(vcc));
defparam \mem[0][5] .is_wysiwyg = "true";
defparam \mem[0][5] .power_up = "low";

dffeas \mem[0][6] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_6_0),
	.prn(vcc));
defparam \mem[0][6] .is_wysiwyg = "true";
defparam \mem[0][6] .power_up = "low";

dffeas \mem[0][7] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_7_0),
	.prn(vcc));
defparam \mem[0][7] .is_wysiwyg = "true";
defparam \mem[0][7] .power_up = "low";

dffeas \mem[0][8] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_8_0),
	.prn(vcc));
defparam \mem[0][8] .is_wysiwyg = "true";
defparam \mem[0][8] .power_up = "low";

dffeas \mem[0][9] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_9_0),
	.prn(vcc));
defparam \mem[0][9] .is_wysiwyg = "true";
defparam \mem[0][9] .power_up = "low";

dffeas \mem[0][10] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_10_0),
	.prn(vcc));
defparam \mem[0][10] .is_wysiwyg = "true";
defparam \mem[0][10] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!h2f_RREADY_0),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem_used[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'h02EA02EA02EA02EA;
defparam \mem_used[1]~1 .shared_arith = "off";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[1]~q ),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~0 (
	.dataa(!h2f_RREADY_0),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem_used[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~0 .extended_lut = "off";
defparam \mem_used[0]~0 .lut_mask = 64'h2B1F2B1F2B1F2B1F;
defparam \mem_used[0]~0 .shared_arith = "off";

dffeas \mem[1][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][0]~q ),
	.prn(vcc));
defparam \mem[1][0] .is_wysiwyg = "true";
defparam \mem[1][0] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!av_readdata_pre_0),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h4747474747474747;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!h2f_RREADY_0),
	.datab(!mem_used_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \always0~0 .shared_arith = "off";

dffeas \mem[1][1] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][1]~q ),
	.prn(vcc));
defparam \mem[1][1] .is_wysiwyg = "true";
defparam \mem[1][1] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!av_readdata_pre_1),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h4747474747474747;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[1][2] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][2]~q ),
	.prn(vcc));
defparam \mem[1][2] .is_wysiwyg = "true";
defparam \mem[1][2] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!av_readdata_pre_2),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h4747474747474747;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[1][3] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][3]~q ),
	.prn(vcc));
defparam \mem[1][3] .is_wysiwyg = "true";
defparam \mem[1][3] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!av_readdata_pre_3),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h4747474747474747;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][4] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][4]~q ),
	.prn(vcc));
defparam \mem[1][4] .is_wysiwyg = "true";
defparam \mem[1][4] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!av_readdata_pre_4),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h4747474747474747;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][5] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][5]~q ),
	.prn(vcc));
defparam \mem[1][5] .is_wysiwyg = "true";
defparam \mem[1][5] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!av_readdata_pre_5),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][5]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h4747474747474747;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][6] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][6]~q ),
	.prn(vcc));
defparam \mem[1][6] .is_wysiwyg = "true";
defparam \mem[1][6] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!av_readdata_pre_6),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][6]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h4747474747474747;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[1][7] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][7]~q ),
	.prn(vcc));
defparam \mem[1][7] .is_wysiwyg = "true";
defparam \mem[1][7] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!av_readdata_pre_7),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h4747474747474747;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[1][8] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][8]~q ),
	.prn(vcc));
defparam \mem[1][8] .is_wysiwyg = "true";
defparam \mem[1][8] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!av_readdata_pre_8),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][8]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h4747474747474747;
defparam \mem~8 .shared_arith = "off";

dffeas \mem[1][9] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][9]~q ),
	.prn(vcc));
defparam \mem[1][9] .is_wysiwyg = "true";
defparam \mem[1][9] .power_up = "low";

cyclonev_lcell_comb \mem~9 (
	.dataa(!av_readdata_pre_9),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][9]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~9 .extended_lut = "off";
defparam \mem~9 .lut_mask = 64'h4747474747474747;
defparam \mem~9 .shared_arith = "off";

dffeas \mem[1][10] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][10]~q ),
	.prn(vcc));
defparam \mem[1][10] .is_wysiwyg = "true";
defparam \mem[1][10] .power_up = "low";

cyclonev_lcell_comb \mem~10 (
	.dataa(!av_readdata_pre_10),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][10]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~10 .extended_lut = "off";
defparam \mem~10 .lut_mask = 64'h4747474747474747;
defparam \mem~10 .shared_arith = "off";

endmodule

module spw_babasu_altera_avalon_sc_fifo_9 (
	h2f_RREADY_0,
	waitrequest_reset_override,
	in_data_reg_69,
	mem_used_1,
	wait_latency_counter_1,
	wait_latency_counter_0,
	out_valid_reg,
	stateST_UNCOMP_WR_SUBBURST,
	empty,
	mem_66_0,
	mem_used_0,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	last_packet_beat,
	mem_130_0,
	mem_105_0,
	mem_106_0,
	mem_107_0,
	mem_108_0,
	mem_109_0,
	mem_110_0,
	mem_111_0,
	mem_112_0,
	mem_113_0,
	mem_114_0,
	mem_115_0,
	mem_116_0,
	reset,
	nxt_out_eop,
	out_byte_cnt_reg_2,
	write,
	write1,
	out_uncomp_byte_cnt_reg_6,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_RREADY_0;
input 	waitrequest_reset_override;
input 	in_data_reg_69;
output 	mem_used_1;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	out_valid_reg;
input 	stateST_UNCOMP_WR_SUBBURST;
input 	empty;
output 	mem_66_0;
output 	mem_used_0;
output 	mem_78_0;
output 	mem_77_0;
output 	mem_76_0;
output 	mem_75_0;
output 	mem_74_0;
input 	last_packet_beat;
output 	mem_130_0;
output 	mem_105_0;
output 	mem_106_0;
output 	mem_107_0;
output 	mem_108_0;
output 	mem_109_0;
output 	mem_110_0;
output 	mem_111_0;
output 	mem_112_0;
output 	mem_113_0;
output 	mem_114_0;
output 	mem_115_0;
output 	mem_116_0;
input 	reset;
input 	nxt_out_eop;
input 	out_byte_cnt_reg_2;
output 	write;
output 	write1;
input 	out_uncomp_byte_cnt_reg_6;
input 	out_uncomp_byte_cnt_reg_5;
input 	out_uncomp_byte_cnt_reg_4;
input 	out_uncomp_byte_cnt_reg_3;
input 	out_uncomp_byte_cnt_reg_2;
input 	in_data_reg_105;
input 	in_data_reg_106;
input 	in_data_reg_107;
input 	in_data_reg_108;
input 	in_data_reg_109;
input 	in_data_reg_110;
input 	in_data_reg_111;
input 	in_data_reg_112;
input 	in_data_reg_113;
input 	in_data_reg_114;
input 	in_data_reg_115;
input 	in_data_reg_116;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read~0_combout ;
wire \mem_used[1]~0_combout ;
wire \mem[1][69]~q ;
wire \mem~0_combout ;
wire \always0~0_combout ;
wire \mem_used[0]~1_combout ;
wire \mem[1][78]~q ;
wire \mem~1_combout ;
wire \mem[1][77]~q ;
wire \mem~2_combout ;
wire \mem[1][76]~q ;
wire \mem~3_combout ;
wire \mem[1][75]~q ;
wire \mem~4_combout ;
wire \mem[1][74]~q ;
wire \mem~5_combout ;
wire \mem[1][130]~q ;
wire \mem~6_combout ;
wire \mem[1][105]~q ;
wire \mem~7_combout ;
wire \mem[1][106]~q ;
wire \mem~8_combout ;
wire \mem[1][107]~q ;
wire \mem~9_combout ;
wire \mem[1][108]~q ;
wire \mem~10_combout ;
wire \mem[1][109]~q ;
wire \mem~11_combout ;
wire \mem[1][110]~q ;
wire \mem~12_combout ;
wire \mem[1][111]~q ;
wire \mem~13_combout ;
wire \mem[1][112]~q ;
wire \mem~14_combout ;
wire \mem[1][113]~q ;
wire \mem~15_combout ;
wire \mem[1][114]~q ;
wire \mem~16_combout ;
wire \mem[1][115]~q ;
wire \mem~17_combout ;
wire \mem[1][116]~q ;
wire \mem~18_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][66] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_66_0),
	.prn(vcc));
defparam \mem[0][66] .is_wysiwyg = "true";
defparam \mem[0][66] .power_up = "low";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][78] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_78_0),
	.prn(vcc));
defparam \mem[0][78] .is_wysiwyg = "true";
defparam \mem[0][78] .power_up = "low";

dffeas \mem[0][77] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_77_0),
	.prn(vcc));
defparam \mem[0][77] .is_wysiwyg = "true";
defparam \mem[0][77] .power_up = "low";

dffeas \mem[0][76] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_76_0),
	.prn(vcc));
defparam \mem[0][76] .is_wysiwyg = "true";
defparam \mem[0][76] .power_up = "low";

dffeas \mem[0][75] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_75_0),
	.prn(vcc));
defparam \mem[0][75] .is_wysiwyg = "true";
defparam \mem[0][75] .power_up = "low";

dffeas \mem[0][74] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_74_0),
	.prn(vcc));
defparam \mem[0][74] .is_wysiwyg = "true";
defparam \mem[0][74] .power_up = "low";

dffeas \mem[0][130] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_130_0),
	.prn(vcc));
defparam \mem[0][130] .is_wysiwyg = "true";
defparam \mem[0][130] .power_up = "low";

dffeas \mem[0][105] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_105_0),
	.prn(vcc));
defparam \mem[0][105] .is_wysiwyg = "true";
defparam \mem[0][105] .power_up = "low";

dffeas \mem[0][106] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_106_0),
	.prn(vcc));
defparam \mem[0][106] .is_wysiwyg = "true";
defparam \mem[0][106] .power_up = "low";

dffeas \mem[0][107] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_107_0),
	.prn(vcc));
defparam \mem[0][107] .is_wysiwyg = "true";
defparam \mem[0][107] .power_up = "low";

dffeas \mem[0][108] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_108_0),
	.prn(vcc));
defparam \mem[0][108] .is_wysiwyg = "true";
defparam \mem[0][108] .power_up = "low";

dffeas \mem[0][109] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_109_0),
	.prn(vcc));
defparam \mem[0][109] .is_wysiwyg = "true";
defparam \mem[0][109] .power_up = "low";

dffeas \mem[0][110] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_110_0),
	.prn(vcc));
defparam \mem[0][110] .is_wysiwyg = "true";
defparam \mem[0][110] .power_up = "low";

dffeas \mem[0][111] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_111_0),
	.prn(vcc));
defparam \mem[0][111] .is_wysiwyg = "true";
defparam \mem[0][111] .power_up = "low";

dffeas \mem[0][112] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_112_0),
	.prn(vcc));
defparam \mem[0][112] .is_wysiwyg = "true";
defparam \mem[0][112] .power_up = "low";

dffeas \mem[0][113] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_113_0),
	.prn(vcc));
defparam \mem[0][113] .is_wysiwyg = "true";
defparam \mem[0][113] .power_up = "low";

dffeas \mem[0][114] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_114_0),
	.prn(vcc));
defparam \mem[0][114] .is_wysiwyg = "true";
defparam \mem[0][114] .power_up = "low";

dffeas \mem[0][115] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_115_0),
	.prn(vcc));
defparam \mem[0][115] .is_wysiwyg = "true";
defparam \mem[0][115] .power_up = "low";

dffeas \mem[0][116] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_116_0),
	.prn(vcc));
defparam \mem[0][116] .is_wysiwyg = "true";
defparam \mem[0][116] .power_up = "low";

cyclonev_lcell_comb \write~0 (
	.dataa(!waitrequest_reset_override),
	.datab(!in_data_reg_69),
	.datac(!mem_used_1),
	.datad(!out_valid_reg),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'h0010001000100010;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \write~1 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!write),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write1),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~1 .extended_lut = "off";
defparam \write~1 .lut_mask = 64'h0202020202020202;
defparam \write~1 .shared_arith = "off";

cyclonev_lcell_comb \read~0 (
	.dataa(!h2f_RREADY_0),
	.datab(!empty),
	.datac(!last_packet_beat),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h4040404040404040;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!\read~0_combout ),
	.datad(!write1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'h5431543154315431;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][69] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][69]~q ),
	.prn(vcc));
defparam \mem[1][69] .is_wysiwyg = "true";
defparam \mem[1][69] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!in_data_reg_69),
	.datab(!mem_used_1),
	.datac(!\mem[1][69]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h4747474747474747;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!mem_used_0),
	.datab(!\read~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!\read~0_combout ),
	.datad(!write1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'h31FF31FF31FF31FF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem[1][78] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][78]~q ),
	.prn(vcc));
defparam \mem[1][78] .is_wysiwyg = "true";
defparam \mem[1][78] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_6),
	.datad(!\mem[1][78]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h0257025702570257;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[1][77] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][77]~q ),
	.prn(vcc));
defparam \mem[1][77] .is_wysiwyg = "true";
defparam \mem[1][77] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\mem[1][77]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h0257025702570257;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[1][76] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][76]~q ),
	.prn(vcc));
defparam \mem[1][76] .is_wysiwyg = "true";
defparam \mem[1][76] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!\mem[1][76]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h0257025702570257;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][75] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][75]~q ),
	.prn(vcc));
defparam \mem[1][75] .is_wysiwyg = "true";
defparam \mem[1][75] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\mem[1][75]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h0257025702570257;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][74] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][74]~q ),
	.prn(vcc));
defparam \mem[1][74] .is_wysiwyg = "true";
defparam \mem[1][74] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_byte_cnt_reg_2),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(!\mem[1][74]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h082A5D7F082A5D7F;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][130] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][130]~q ),
	.prn(vcc));
defparam \mem[1][130] .is_wysiwyg = "true";
defparam \mem[1][130] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!mem_used_1),
	.datab(!nxt_out_eop),
	.datac(!\mem[1][130]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h2727272727272727;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[1][105] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][105]~q ),
	.prn(vcc));
defparam \mem[1][105] .is_wysiwyg = "true";
defparam \mem[1][105] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][105]~q ),
	.datac(!in_data_reg_105),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[1][106] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][106]~q ),
	.prn(vcc));
defparam \mem[1][106] .is_wysiwyg = "true";
defparam \mem[1][106] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][106]~q ),
	.datac(!in_data_reg_106),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~8 .shared_arith = "off";

dffeas \mem[1][107] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][107]~q ),
	.prn(vcc));
defparam \mem[1][107] .is_wysiwyg = "true";
defparam \mem[1][107] .power_up = "low";

cyclonev_lcell_comb \mem~9 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][107]~q ),
	.datac(!in_data_reg_107),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~9 .extended_lut = "off";
defparam \mem~9 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~9 .shared_arith = "off";

dffeas \mem[1][108] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][108]~q ),
	.prn(vcc));
defparam \mem[1][108] .is_wysiwyg = "true";
defparam \mem[1][108] .power_up = "low";

cyclonev_lcell_comb \mem~10 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][108]~q ),
	.datac(!in_data_reg_108),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~10 .extended_lut = "off";
defparam \mem~10 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~10 .shared_arith = "off";

dffeas \mem[1][109] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][109]~q ),
	.prn(vcc));
defparam \mem[1][109] .is_wysiwyg = "true";
defparam \mem[1][109] .power_up = "low";

cyclonev_lcell_comb \mem~11 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][109]~q ),
	.datac(!in_data_reg_109),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~11 .extended_lut = "off";
defparam \mem~11 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~11 .shared_arith = "off";

dffeas \mem[1][110] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][110]~q ),
	.prn(vcc));
defparam \mem[1][110] .is_wysiwyg = "true";
defparam \mem[1][110] .power_up = "low";

cyclonev_lcell_comb \mem~12 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][110]~q ),
	.datac(!in_data_reg_110),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~12 .extended_lut = "off";
defparam \mem~12 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~12 .shared_arith = "off";

dffeas \mem[1][111] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][111]~q ),
	.prn(vcc));
defparam \mem[1][111] .is_wysiwyg = "true";
defparam \mem[1][111] .power_up = "low";

cyclonev_lcell_comb \mem~13 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][111]~q ),
	.datac(!in_data_reg_111),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~13 .extended_lut = "off";
defparam \mem~13 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~13 .shared_arith = "off";

dffeas \mem[1][112] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][112]~q ),
	.prn(vcc));
defparam \mem[1][112] .is_wysiwyg = "true";
defparam \mem[1][112] .power_up = "low";

cyclonev_lcell_comb \mem~14 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][112]~q ),
	.datac(!in_data_reg_112),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~14 .extended_lut = "off";
defparam \mem~14 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~14 .shared_arith = "off";

dffeas \mem[1][113] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][113]~q ),
	.prn(vcc));
defparam \mem[1][113] .is_wysiwyg = "true";
defparam \mem[1][113] .power_up = "low";

cyclonev_lcell_comb \mem~15 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][113]~q ),
	.datac(!in_data_reg_113),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~15 .extended_lut = "off";
defparam \mem~15 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~15 .shared_arith = "off";

dffeas \mem[1][114] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][114]~q ),
	.prn(vcc));
defparam \mem[1][114] .is_wysiwyg = "true";
defparam \mem[1][114] .power_up = "low";

cyclonev_lcell_comb \mem~16 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][114]~q ),
	.datac(!in_data_reg_114),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~16 .extended_lut = "off";
defparam \mem~16 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~16 .shared_arith = "off";

dffeas \mem[1][115] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][115]~q ),
	.prn(vcc));
defparam \mem[1][115] .is_wysiwyg = "true";
defparam \mem[1][115] .power_up = "low";

cyclonev_lcell_comb \mem~17 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][115]~q ),
	.datac(!in_data_reg_115),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~17 .extended_lut = "off";
defparam \mem~17 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~17 .shared_arith = "off";

dffeas \mem[1][116] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][116]~q ),
	.prn(vcc));
defparam \mem[1][116] .is_wysiwyg = "true";
defparam \mem[1][116] .power_up = "low";

cyclonev_lcell_comb \mem~18 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][116]~q ),
	.datac(!in_data_reg_116),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~18 .extended_lut = "off";
defparam \mem~18 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~18 .shared_arith = "off";

endmodule

module spw_babasu_altera_avalon_sc_fifo_10 (
	read_latency_shift_reg_0,
	mem_used_0,
	mem_129_0,
	mem_used_01,
	av_readdata_pre_0,
	mem_0_0,
	reset,
	WideOr0,
	clk)/* synthesis synthesis_greybox=0 */;
input 	read_latency_shift_reg_0;
output 	mem_used_0;
input 	mem_129_0;
input 	mem_used_01;
input 	av_readdata_pre_0;
output 	mem_0_0;
input 	reset;
input 	WideOr0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~q ;
wire \mem_used[0]~0_combout ;
wire \mem[1][0]~q ;
wire \mem~0_combout ;
wire \mem[0][0]~1_combout ;


dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][0] (
	.clk(clk),
	.d(\mem[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_0_0),
	.prn(vcc));
defparam \mem[0][0] .is_wysiwyg = "true";
defparam \mem[0][0] .power_up = "low";

cyclonev_lcell_comb \read~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_129_0),
	.datad(!mem_used_01),
	.datae(!WideOr0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h0000777000007770;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!\mem_used[1]~q ),
	.datad(!\read~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'h1F001F001F001F00;
defparam \mem_used[1]~1 .shared_arith = "off";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[1]~q ),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!\mem_used[1]~q ),
	.datad(!\read~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~0 .extended_lut = "off";
defparam \mem_used[0]~0 .lut_mask = 64'h731F731F731F731F;
defparam \mem_used[0]~0 .shared_arith = "off";

dffeas \mem[1][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][0]~q ),
	.prn(vcc));
defparam \mem[1][0] .is_wysiwyg = "true";
defparam \mem[1][0] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!av_readdata_pre_0),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h4747474747474747;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \mem[0][0]~1 (
	.dataa(!mem_used_0),
	.datab(!mem_0_0),
	.datac(!\read~0_combout ),
	.datad(!\mem~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem[0][0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem[0][0]~1 .extended_lut = "off";
defparam \mem[0][0]~1 .lut_mask = 64'h10BF10BF10BF10BF;
defparam \mem[0][0]~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_avalon_sc_fifo_11 (
	out_valid_reg,
	mem_used_1,
	WideOr0,
	in_data_reg_68,
	stateST_UNCOMP_WR_SUBBURST,
	mem_129_0,
	mem_used_0,
	mem_68_0,
	mem_66_0,
	comb,
	mem_130_0,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	mem_105_0,
	mem_106_0,
	mem_107_0,
	mem_108_0,
	mem_109_0,
	mem_110_0,
	mem_111_0,
	mem_112_0,
	mem_113_0,
	mem_114_0,
	mem_115_0,
	mem_116_0,
	reset,
	nxt_out_eop,
	last_packet_beat,
	WideOr01,
	read,
	cp_ready,
	in_data_reg_69,
	rf_source_valid,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_6,
	sink_ready,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	clk)/* synthesis synthesis_greybox=0 */;
input 	out_valid_reg;
output 	mem_used_1;
input 	WideOr0;
input 	in_data_reg_68;
input 	stateST_UNCOMP_WR_SUBBURST;
output 	mem_129_0;
output 	mem_used_0;
output 	mem_68_0;
output 	mem_66_0;
input 	comb;
output 	mem_130_0;
output 	mem_78_0;
output 	mem_77_0;
output 	mem_76_0;
output 	mem_75_0;
output 	mem_74_0;
output 	mem_105_0;
output 	mem_106_0;
output 	mem_107_0;
output 	mem_108_0;
output 	mem_109_0;
output 	mem_110_0;
output 	mem_111_0;
output 	mem_112_0;
output 	mem_113_0;
output 	mem_114_0;
output 	mem_115_0;
output 	mem_116_0;
input 	reset;
input 	nxt_out_eop;
input 	last_packet_beat;
input 	WideOr01;
output 	read;
input 	cp_ready;
input 	in_data_reg_69;
input 	rf_source_valid;
input 	out_byte_cnt_reg_2;
input 	out_uncomp_byte_cnt_reg_3;
input 	out_uncomp_byte_cnt_reg_2;
input 	out_uncomp_byte_cnt_reg_4;
input 	out_uncomp_byte_cnt_reg_5;
input 	out_uncomp_byte_cnt_reg_6;
input 	sink_ready;
input 	in_data_reg_105;
input 	in_data_reg_106;
input 	in_data_reg_107;
input 	in_data_reg_108;
input 	in_data_reg_109;
input 	in_data_reg_110;
input 	in_data_reg_111;
input 	in_data_reg_112;
input 	in_data_reg_113;
input 	in_data_reg_114;
input 	in_data_reg_115;
input 	in_data_reg_116;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \write~0_combout ;
wire \mem_used[1]~0_combout ;
wire \mem[1][129]~q ;
wire \mem~20_combout ;
wire \always0~0_combout ;
wire \mem_used[0]~1_combout ;
wire \mem[1][68]~q ;
wire \mem~0_combout ;
wire \mem[1][69]~q ;
wire \mem~1_combout ;
wire \mem[1][130]~q ;
wire \mem~2_combout ;
wire \mem[1][78]~q ;
wire \mem~3_combout ;
wire \mem[1][77]~q ;
wire \mem~4_combout ;
wire \mem[1][76]~q ;
wire \mem~5_combout ;
wire \mem[1][75]~q ;
wire \mem~6_combout ;
wire \mem[1][74]~q ;
wire \mem~7_combout ;
wire \mem[1][105]~q ;
wire \mem~8_combout ;
wire \mem[1][106]~q ;
wire \mem~9_combout ;
wire \mem[1][107]~q ;
wire \mem~10_combout ;
wire \mem[1][108]~q ;
wire \mem~11_combout ;
wire \mem[1][109]~q ;
wire \mem~12_combout ;
wire \mem[1][110]~q ;
wire \mem~13_combout ;
wire \mem[1][111]~q ;
wire \mem~14_combout ;
wire \mem[1][112]~q ;
wire \mem~15_combout ;
wire \mem[1][113]~q ;
wire \mem~16_combout ;
wire \mem[1][114]~q ;
wire \mem~17_combout ;
wire \mem[1][115]~q ;
wire \mem~18_combout ;
wire \mem[1][116]~q ;
wire \mem~19_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][129] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_129_0),
	.prn(vcc));
defparam \mem[0][129] .is_wysiwyg = "true";
defparam \mem[0][129] .power_up = "low";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][68] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_68_0),
	.prn(vcc));
defparam \mem[0][68] .is_wysiwyg = "true";
defparam \mem[0][68] .power_up = "low";

dffeas \mem[0][66] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_66_0),
	.prn(vcc));
defparam \mem[0][66] .is_wysiwyg = "true";
defparam \mem[0][66] .power_up = "low";

dffeas \mem[0][130] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_130_0),
	.prn(vcc));
defparam \mem[0][130] .is_wysiwyg = "true";
defparam \mem[0][130] .power_up = "low";

dffeas \mem[0][78] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_78_0),
	.prn(vcc));
defparam \mem[0][78] .is_wysiwyg = "true";
defparam \mem[0][78] .power_up = "low";

dffeas \mem[0][77] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_77_0),
	.prn(vcc));
defparam \mem[0][77] .is_wysiwyg = "true";
defparam \mem[0][77] .power_up = "low";

dffeas \mem[0][76] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_76_0),
	.prn(vcc));
defparam \mem[0][76] .is_wysiwyg = "true";
defparam \mem[0][76] .power_up = "low";

dffeas \mem[0][75] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_75_0),
	.prn(vcc));
defparam \mem[0][75] .is_wysiwyg = "true";
defparam \mem[0][75] .power_up = "low";

dffeas \mem[0][74] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_74_0),
	.prn(vcc));
defparam \mem[0][74] .is_wysiwyg = "true";
defparam \mem[0][74] .power_up = "low";

dffeas \mem[0][105] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_105_0),
	.prn(vcc));
defparam \mem[0][105] .is_wysiwyg = "true";
defparam \mem[0][105] .power_up = "low";

dffeas \mem[0][106] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_106_0),
	.prn(vcc));
defparam \mem[0][106] .is_wysiwyg = "true";
defparam \mem[0][106] .power_up = "low";

dffeas \mem[0][107] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_107_0),
	.prn(vcc));
defparam \mem[0][107] .is_wysiwyg = "true";
defparam \mem[0][107] .power_up = "low";

dffeas \mem[0][108] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_108_0),
	.prn(vcc));
defparam \mem[0][108] .is_wysiwyg = "true";
defparam \mem[0][108] .power_up = "low";

dffeas \mem[0][109] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_109_0),
	.prn(vcc));
defparam \mem[0][109] .is_wysiwyg = "true";
defparam \mem[0][109] .power_up = "low";

dffeas \mem[0][110] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_110_0),
	.prn(vcc));
defparam \mem[0][110] .is_wysiwyg = "true";
defparam \mem[0][110] .power_up = "low";

dffeas \mem[0][111] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_111_0),
	.prn(vcc));
defparam \mem[0][111] .is_wysiwyg = "true";
defparam \mem[0][111] .power_up = "low";

dffeas \mem[0][112] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_112_0),
	.prn(vcc));
defparam \mem[0][112] .is_wysiwyg = "true";
defparam \mem[0][112] .power_up = "low";

dffeas \mem[0][113] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_113_0),
	.prn(vcc));
defparam \mem[0][113] .is_wysiwyg = "true";
defparam \mem[0][113] .power_up = "low";

dffeas \mem[0][114] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_114_0),
	.prn(vcc));
defparam \mem[0][114] .is_wysiwyg = "true";
defparam \mem[0][114] .power_up = "low";

dffeas \mem[0][115] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_115_0),
	.prn(vcc));
defparam \mem[0][115] .is_wysiwyg = "true";
defparam \mem[0][115] .power_up = "low";

dffeas \mem[0][116] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_116_0),
	.prn(vcc));
defparam \mem[0][116] .is_wysiwyg = "true";
defparam \mem[0][116] .power_up = "low";

cyclonev_lcell_comb \read~0 (
	.dataa(!comb),
	.datab(!WideOr01),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h1111111111111111;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \write~0 (
	.dataa(!mem_used_1),
	.datab(!WideOr0),
	.datac(!cp_ready),
	.datad(!rf_source_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'h008A008A008A008A;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!last_packet_beat),
	.datad(!read),
	.datae(!\write~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'h5505335355053353;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][129] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][129]~q ),
	.prn(vcc));
defparam \mem[1][129] .is_wysiwyg = "true";
defparam \mem[1][129] .power_up = "low";

cyclonev_lcell_comb \mem~20 (
	.dataa(!WideOr0),
	.datab(!out_valid_reg),
	.datac(!\mem[1][129]~q ),
	.datad(!in_data_reg_68),
	.datae(!mem_used_1),
	.dataf(!nxt_out_eop),
	.datag(!in_data_reg_69),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~20 .extended_lut = "on";
defparam \mem~20 .lut_mask = 64'h02020F0F02330F0F;
defparam \mem~20 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!mem_used_0),
	.datab(!sink_ready),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!\write~0_combout ),
	.datad(!sink_ready),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'h3F1F3F1F3F1F3F1F;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem[1][68] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][68]~q ),
	.prn(vcc));
defparam \mem[1][68] .is_wysiwyg = "true";
defparam \mem[1][68] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!mem_used_1),
	.datab(!in_data_reg_68),
	.datac(!\mem[1][68]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h2727272727272727;
defparam \mem~0 .shared_arith = "off";

dffeas \mem[1][69] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][69]~q ),
	.prn(vcc));
defparam \mem[1][69] .is_wysiwyg = "true";
defparam \mem[1][69] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!mem_used_1),
	.datab(!in_data_reg_69),
	.datac(!\mem[1][69]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h2727272727272727;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[1][130] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][130]~q ),
	.prn(vcc));
defparam \mem[1][130] .is_wysiwyg = "true";
defparam \mem[1][130] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!mem_used_1),
	.datab(!nxt_out_eop),
	.datac(!\mem[1][130]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h2727272727272727;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[1][78] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][78]~q ),
	.prn(vcc));
defparam \mem[1][78] .is_wysiwyg = "true";
defparam \mem[1][78] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_6),
	.datad(!\mem[1][78]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h0257025702570257;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][77] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][77]~q ),
	.prn(vcc));
defparam \mem[1][77] .is_wysiwyg = "true";
defparam \mem[1][77] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\mem[1][77]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h0257025702570257;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][76] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][76]~q ),
	.prn(vcc));
defparam \mem[1][76] .is_wysiwyg = "true";
defparam \mem[1][76] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!\mem[1][76]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h0257025702570257;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][75] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][75]~q ),
	.prn(vcc));
defparam \mem[1][75] .is_wysiwyg = "true";
defparam \mem[1][75] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\mem[1][75]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h0257025702570257;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[1][74] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][74]~q ),
	.prn(vcc));
defparam \mem[1][74] .is_wysiwyg = "true";
defparam \mem[1][74] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_byte_cnt_reg_2),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(!\mem[1][74]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h082A5D7F082A5D7F;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[1][105] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][105]~q ),
	.prn(vcc));
defparam \mem[1][105] .is_wysiwyg = "true";
defparam \mem[1][105] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][105]~q ),
	.datac(!in_data_reg_105),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~8 .shared_arith = "off";

dffeas \mem[1][106] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][106]~q ),
	.prn(vcc));
defparam \mem[1][106] .is_wysiwyg = "true";
defparam \mem[1][106] .power_up = "low";

cyclonev_lcell_comb \mem~9 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][106]~q ),
	.datac(!in_data_reg_106),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~9 .extended_lut = "off";
defparam \mem~9 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~9 .shared_arith = "off";

dffeas \mem[1][107] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][107]~q ),
	.prn(vcc));
defparam \mem[1][107] .is_wysiwyg = "true";
defparam \mem[1][107] .power_up = "low";

cyclonev_lcell_comb \mem~10 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][107]~q ),
	.datac(!in_data_reg_107),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~10 .extended_lut = "off";
defparam \mem~10 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~10 .shared_arith = "off";

dffeas \mem[1][108] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][108]~q ),
	.prn(vcc));
defparam \mem[1][108] .is_wysiwyg = "true";
defparam \mem[1][108] .power_up = "low";

cyclonev_lcell_comb \mem~11 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][108]~q ),
	.datac(!in_data_reg_108),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~11 .extended_lut = "off";
defparam \mem~11 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~11 .shared_arith = "off";

dffeas \mem[1][109] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][109]~q ),
	.prn(vcc));
defparam \mem[1][109] .is_wysiwyg = "true";
defparam \mem[1][109] .power_up = "low";

cyclonev_lcell_comb \mem~12 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][109]~q ),
	.datac(!in_data_reg_109),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~12 .extended_lut = "off";
defparam \mem~12 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~12 .shared_arith = "off";

dffeas \mem[1][110] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][110]~q ),
	.prn(vcc));
defparam \mem[1][110] .is_wysiwyg = "true";
defparam \mem[1][110] .power_up = "low";

cyclonev_lcell_comb \mem~13 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][110]~q ),
	.datac(!in_data_reg_110),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~13 .extended_lut = "off";
defparam \mem~13 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~13 .shared_arith = "off";

dffeas \mem[1][111] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][111]~q ),
	.prn(vcc));
defparam \mem[1][111] .is_wysiwyg = "true";
defparam \mem[1][111] .power_up = "low";

cyclonev_lcell_comb \mem~14 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][111]~q ),
	.datac(!in_data_reg_111),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~14 .extended_lut = "off";
defparam \mem~14 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~14 .shared_arith = "off";

dffeas \mem[1][112] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][112]~q ),
	.prn(vcc));
defparam \mem[1][112] .is_wysiwyg = "true";
defparam \mem[1][112] .power_up = "low";

cyclonev_lcell_comb \mem~15 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][112]~q ),
	.datac(!in_data_reg_112),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~15 .extended_lut = "off";
defparam \mem~15 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~15 .shared_arith = "off";

dffeas \mem[1][113] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][113]~q ),
	.prn(vcc));
defparam \mem[1][113] .is_wysiwyg = "true";
defparam \mem[1][113] .power_up = "low";

cyclonev_lcell_comb \mem~16 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][113]~q ),
	.datac(!in_data_reg_113),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~16 .extended_lut = "off";
defparam \mem~16 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~16 .shared_arith = "off";

dffeas \mem[1][114] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][114]~q ),
	.prn(vcc));
defparam \mem[1][114] .is_wysiwyg = "true";
defparam \mem[1][114] .power_up = "low";

cyclonev_lcell_comb \mem~17 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][114]~q ),
	.datac(!in_data_reg_114),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~17 .extended_lut = "off";
defparam \mem~17 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~17 .shared_arith = "off";

dffeas \mem[1][115] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][115]~q ),
	.prn(vcc));
defparam \mem[1][115] .is_wysiwyg = "true";
defparam \mem[1][115] .power_up = "low";

cyclonev_lcell_comb \mem~18 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][115]~q ),
	.datac(!in_data_reg_115),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~18 .extended_lut = "off";
defparam \mem~18 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~18 .shared_arith = "off";

dffeas \mem[1][116] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][116]~q ),
	.prn(vcc));
defparam \mem[1][116] .is_wysiwyg = "true";
defparam \mem[1][116] .power_up = "low";

cyclonev_lcell_comb \mem~19 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][116]~q ),
	.datac(!in_data_reg_116),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~19 .extended_lut = "off";
defparam \mem~19 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~19 .shared_arith = "off";

endmodule

module spw_babasu_altera_avalon_sc_fifo_12 (
	read_latency_shift_reg_0,
	mem_used_0,
	mem_129_0,
	mem_used_01,
	av_readdata_pre_0,
	mem_0_0,
	reset,
	WideOr0,
	clk)/* synthesis synthesis_greybox=0 */;
input 	read_latency_shift_reg_0;
output 	mem_used_0;
input 	mem_129_0;
input 	mem_used_01;
input 	av_readdata_pre_0;
output 	mem_0_0;
input 	reset;
input 	WideOr0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~q ;
wire \mem_used[0]~0_combout ;
wire \mem[1][0]~q ;
wire \mem~0_combout ;
wire \mem[0][0]~1_combout ;


dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][0] (
	.clk(clk),
	.d(\mem[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_0_0),
	.prn(vcc));
defparam \mem[0][0] .is_wysiwyg = "true";
defparam \mem[0][0] .power_up = "low";

cyclonev_lcell_comb \read~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_129_0),
	.datad(!mem_used_01),
	.datae(!WideOr0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h0000777000007770;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!\mem_used[1]~q ),
	.datad(!\read~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'h1F001F001F001F00;
defparam \mem_used[1]~1 .shared_arith = "off";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[1]~q ),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!\mem_used[1]~q ),
	.datad(!\read~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~0 .extended_lut = "off";
defparam \mem_used[0]~0 .lut_mask = 64'h731F731F731F731F;
defparam \mem_used[0]~0 .shared_arith = "off";

dffeas \mem[1][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][0]~q ),
	.prn(vcc));
defparam \mem[1][0] .is_wysiwyg = "true";
defparam \mem[1][0] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!av_readdata_pre_0),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h4747474747474747;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \mem[0][0]~1 (
	.dataa(!mem_used_0),
	.datab(!mem_0_0),
	.datac(!\read~0_combout ),
	.datad(!\mem~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem[0][0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem[0][0]~1 .extended_lut = "off";
defparam \mem[0][0]~1 .lut_mask = 64'h10BF10BF10BF10BF;
defparam \mem[0][0]~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_avalon_sc_fifo_13 (
	out_valid_reg,
	mem_used_1,
	WideOr0,
	in_data_reg_68,
	stateST_UNCOMP_WR_SUBBURST,
	mem_129_0,
	mem_used_0,
	mem_68_0,
	mem_66_0,
	comb,
	mem_130_0,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	mem_105_0,
	mem_106_0,
	mem_107_0,
	mem_108_0,
	mem_109_0,
	mem_110_0,
	mem_111_0,
	mem_112_0,
	mem_113_0,
	mem_114_0,
	mem_115_0,
	mem_116_0,
	reset,
	nxt_out_eop,
	last_packet_beat,
	WideOr01,
	read,
	cp_ready,
	in_data_reg_69,
	rf_source_valid,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_6,
	sink_ready,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	clk)/* synthesis synthesis_greybox=0 */;
input 	out_valid_reg;
output 	mem_used_1;
input 	WideOr0;
input 	in_data_reg_68;
input 	stateST_UNCOMP_WR_SUBBURST;
output 	mem_129_0;
output 	mem_used_0;
output 	mem_68_0;
output 	mem_66_0;
input 	comb;
output 	mem_130_0;
output 	mem_78_0;
output 	mem_77_0;
output 	mem_76_0;
output 	mem_75_0;
output 	mem_74_0;
output 	mem_105_0;
output 	mem_106_0;
output 	mem_107_0;
output 	mem_108_0;
output 	mem_109_0;
output 	mem_110_0;
output 	mem_111_0;
output 	mem_112_0;
output 	mem_113_0;
output 	mem_114_0;
output 	mem_115_0;
output 	mem_116_0;
input 	reset;
input 	nxt_out_eop;
input 	last_packet_beat;
input 	WideOr01;
output 	read;
input 	cp_ready;
input 	in_data_reg_69;
input 	rf_source_valid;
input 	out_byte_cnt_reg_2;
input 	out_uncomp_byte_cnt_reg_3;
input 	out_uncomp_byte_cnt_reg_2;
input 	out_uncomp_byte_cnt_reg_4;
input 	out_uncomp_byte_cnt_reg_5;
input 	out_uncomp_byte_cnt_reg_6;
input 	sink_ready;
input 	in_data_reg_105;
input 	in_data_reg_106;
input 	in_data_reg_107;
input 	in_data_reg_108;
input 	in_data_reg_109;
input 	in_data_reg_110;
input 	in_data_reg_111;
input 	in_data_reg_112;
input 	in_data_reg_113;
input 	in_data_reg_114;
input 	in_data_reg_115;
input 	in_data_reg_116;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \write~0_combout ;
wire \mem_used[1]~0_combout ;
wire \mem[1][129]~q ;
wire \mem~20_combout ;
wire \always0~0_combout ;
wire \mem_used[0]~1_combout ;
wire \mem[1][68]~q ;
wire \mem~0_combout ;
wire \mem[1][69]~q ;
wire \mem~1_combout ;
wire \mem[1][130]~q ;
wire \mem~2_combout ;
wire \mem[1][78]~q ;
wire \mem~3_combout ;
wire \mem[1][77]~q ;
wire \mem~4_combout ;
wire \mem[1][76]~q ;
wire \mem~5_combout ;
wire \mem[1][75]~q ;
wire \mem~6_combout ;
wire \mem[1][74]~q ;
wire \mem~7_combout ;
wire \mem[1][105]~q ;
wire \mem~8_combout ;
wire \mem[1][106]~q ;
wire \mem~9_combout ;
wire \mem[1][107]~q ;
wire \mem~10_combout ;
wire \mem[1][108]~q ;
wire \mem~11_combout ;
wire \mem[1][109]~q ;
wire \mem~12_combout ;
wire \mem[1][110]~q ;
wire \mem~13_combout ;
wire \mem[1][111]~q ;
wire \mem~14_combout ;
wire \mem[1][112]~q ;
wire \mem~15_combout ;
wire \mem[1][113]~q ;
wire \mem~16_combout ;
wire \mem[1][114]~q ;
wire \mem~17_combout ;
wire \mem[1][115]~q ;
wire \mem~18_combout ;
wire \mem[1][116]~q ;
wire \mem~19_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][129] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_129_0),
	.prn(vcc));
defparam \mem[0][129] .is_wysiwyg = "true";
defparam \mem[0][129] .power_up = "low";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][68] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_68_0),
	.prn(vcc));
defparam \mem[0][68] .is_wysiwyg = "true";
defparam \mem[0][68] .power_up = "low";

dffeas \mem[0][66] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_66_0),
	.prn(vcc));
defparam \mem[0][66] .is_wysiwyg = "true";
defparam \mem[0][66] .power_up = "low";

dffeas \mem[0][130] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_130_0),
	.prn(vcc));
defparam \mem[0][130] .is_wysiwyg = "true";
defparam \mem[0][130] .power_up = "low";

dffeas \mem[0][78] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_78_0),
	.prn(vcc));
defparam \mem[0][78] .is_wysiwyg = "true";
defparam \mem[0][78] .power_up = "low";

dffeas \mem[0][77] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_77_0),
	.prn(vcc));
defparam \mem[0][77] .is_wysiwyg = "true";
defparam \mem[0][77] .power_up = "low";

dffeas \mem[0][76] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_76_0),
	.prn(vcc));
defparam \mem[0][76] .is_wysiwyg = "true";
defparam \mem[0][76] .power_up = "low";

dffeas \mem[0][75] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_75_0),
	.prn(vcc));
defparam \mem[0][75] .is_wysiwyg = "true";
defparam \mem[0][75] .power_up = "low";

dffeas \mem[0][74] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_74_0),
	.prn(vcc));
defparam \mem[0][74] .is_wysiwyg = "true";
defparam \mem[0][74] .power_up = "low";

dffeas \mem[0][105] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_105_0),
	.prn(vcc));
defparam \mem[0][105] .is_wysiwyg = "true";
defparam \mem[0][105] .power_up = "low";

dffeas \mem[0][106] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_106_0),
	.prn(vcc));
defparam \mem[0][106] .is_wysiwyg = "true";
defparam \mem[0][106] .power_up = "low";

dffeas \mem[0][107] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_107_0),
	.prn(vcc));
defparam \mem[0][107] .is_wysiwyg = "true";
defparam \mem[0][107] .power_up = "low";

dffeas \mem[0][108] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_108_0),
	.prn(vcc));
defparam \mem[0][108] .is_wysiwyg = "true";
defparam \mem[0][108] .power_up = "low";

dffeas \mem[0][109] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_109_0),
	.prn(vcc));
defparam \mem[0][109] .is_wysiwyg = "true";
defparam \mem[0][109] .power_up = "low";

dffeas \mem[0][110] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_110_0),
	.prn(vcc));
defparam \mem[0][110] .is_wysiwyg = "true";
defparam \mem[0][110] .power_up = "low";

dffeas \mem[0][111] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_111_0),
	.prn(vcc));
defparam \mem[0][111] .is_wysiwyg = "true";
defparam \mem[0][111] .power_up = "low";

dffeas \mem[0][112] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_112_0),
	.prn(vcc));
defparam \mem[0][112] .is_wysiwyg = "true";
defparam \mem[0][112] .power_up = "low";

dffeas \mem[0][113] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_113_0),
	.prn(vcc));
defparam \mem[0][113] .is_wysiwyg = "true";
defparam \mem[0][113] .power_up = "low";

dffeas \mem[0][114] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_114_0),
	.prn(vcc));
defparam \mem[0][114] .is_wysiwyg = "true";
defparam \mem[0][114] .power_up = "low";

dffeas \mem[0][115] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_115_0),
	.prn(vcc));
defparam \mem[0][115] .is_wysiwyg = "true";
defparam \mem[0][115] .power_up = "low";

dffeas \mem[0][116] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_116_0),
	.prn(vcc));
defparam \mem[0][116] .is_wysiwyg = "true";
defparam \mem[0][116] .power_up = "low";

cyclonev_lcell_comb \read~0 (
	.dataa(!comb),
	.datab(!WideOr01),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h1111111111111111;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \write~0 (
	.dataa(!mem_used_1),
	.datab(!WideOr0),
	.datac(!cp_ready),
	.datad(!rf_source_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'h008A008A008A008A;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!last_packet_beat),
	.datad(!read),
	.datae(!\write~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'h5505335355053353;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][129] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][129]~q ),
	.prn(vcc));
defparam \mem[1][129] .is_wysiwyg = "true";
defparam \mem[1][129] .power_up = "low";

cyclonev_lcell_comb \mem~20 (
	.dataa(!WideOr0),
	.datab(!out_valid_reg),
	.datac(!\mem[1][129]~q ),
	.datad(!in_data_reg_68),
	.datae(!mem_used_1),
	.dataf(!nxt_out_eop),
	.datag(!in_data_reg_69),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~20 .extended_lut = "on";
defparam \mem~20 .lut_mask = 64'h02020F0F02330F0F;
defparam \mem~20 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!mem_used_0),
	.datab(!sink_ready),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!\write~0_combout ),
	.datad(!sink_ready),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'h3F1F3F1F3F1F3F1F;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem[1][68] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][68]~q ),
	.prn(vcc));
defparam \mem[1][68] .is_wysiwyg = "true";
defparam \mem[1][68] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!mem_used_1),
	.datab(!in_data_reg_68),
	.datac(!\mem[1][68]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h2727272727272727;
defparam \mem~0 .shared_arith = "off";

dffeas \mem[1][69] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][69]~q ),
	.prn(vcc));
defparam \mem[1][69] .is_wysiwyg = "true";
defparam \mem[1][69] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!mem_used_1),
	.datab(!in_data_reg_69),
	.datac(!\mem[1][69]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h2727272727272727;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[1][130] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][130]~q ),
	.prn(vcc));
defparam \mem[1][130] .is_wysiwyg = "true";
defparam \mem[1][130] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!mem_used_1),
	.datab(!nxt_out_eop),
	.datac(!\mem[1][130]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h2727272727272727;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[1][78] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][78]~q ),
	.prn(vcc));
defparam \mem[1][78] .is_wysiwyg = "true";
defparam \mem[1][78] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_6),
	.datad(!\mem[1][78]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h0257025702570257;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][77] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][77]~q ),
	.prn(vcc));
defparam \mem[1][77] .is_wysiwyg = "true";
defparam \mem[1][77] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\mem[1][77]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h0257025702570257;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][76] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][76]~q ),
	.prn(vcc));
defparam \mem[1][76] .is_wysiwyg = "true";
defparam \mem[1][76] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!\mem[1][76]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h0257025702570257;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][75] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][75]~q ),
	.prn(vcc));
defparam \mem[1][75] .is_wysiwyg = "true";
defparam \mem[1][75] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\mem[1][75]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h0257025702570257;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[1][74] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][74]~q ),
	.prn(vcc));
defparam \mem[1][74] .is_wysiwyg = "true";
defparam \mem[1][74] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_byte_cnt_reg_2),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(!\mem[1][74]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h082A5D7F082A5D7F;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[1][105] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][105]~q ),
	.prn(vcc));
defparam \mem[1][105] .is_wysiwyg = "true";
defparam \mem[1][105] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][105]~q ),
	.datac(!in_data_reg_105),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~8 .shared_arith = "off";

dffeas \mem[1][106] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][106]~q ),
	.prn(vcc));
defparam \mem[1][106] .is_wysiwyg = "true";
defparam \mem[1][106] .power_up = "low";

cyclonev_lcell_comb \mem~9 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][106]~q ),
	.datac(!in_data_reg_106),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~9 .extended_lut = "off";
defparam \mem~9 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~9 .shared_arith = "off";

dffeas \mem[1][107] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][107]~q ),
	.prn(vcc));
defparam \mem[1][107] .is_wysiwyg = "true";
defparam \mem[1][107] .power_up = "low";

cyclonev_lcell_comb \mem~10 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][107]~q ),
	.datac(!in_data_reg_107),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~10 .extended_lut = "off";
defparam \mem~10 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~10 .shared_arith = "off";

dffeas \mem[1][108] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][108]~q ),
	.prn(vcc));
defparam \mem[1][108] .is_wysiwyg = "true";
defparam \mem[1][108] .power_up = "low";

cyclonev_lcell_comb \mem~11 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][108]~q ),
	.datac(!in_data_reg_108),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~11 .extended_lut = "off";
defparam \mem~11 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~11 .shared_arith = "off";

dffeas \mem[1][109] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][109]~q ),
	.prn(vcc));
defparam \mem[1][109] .is_wysiwyg = "true";
defparam \mem[1][109] .power_up = "low";

cyclonev_lcell_comb \mem~12 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][109]~q ),
	.datac(!in_data_reg_109),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~12 .extended_lut = "off";
defparam \mem~12 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~12 .shared_arith = "off";

dffeas \mem[1][110] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][110]~q ),
	.prn(vcc));
defparam \mem[1][110] .is_wysiwyg = "true";
defparam \mem[1][110] .power_up = "low";

cyclonev_lcell_comb \mem~13 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][110]~q ),
	.datac(!in_data_reg_110),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~13 .extended_lut = "off";
defparam \mem~13 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~13 .shared_arith = "off";

dffeas \mem[1][111] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][111]~q ),
	.prn(vcc));
defparam \mem[1][111] .is_wysiwyg = "true";
defparam \mem[1][111] .power_up = "low";

cyclonev_lcell_comb \mem~14 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][111]~q ),
	.datac(!in_data_reg_111),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~14 .extended_lut = "off";
defparam \mem~14 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~14 .shared_arith = "off";

dffeas \mem[1][112] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][112]~q ),
	.prn(vcc));
defparam \mem[1][112] .is_wysiwyg = "true";
defparam \mem[1][112] .power_up = "low";

cyclonev_lcell_comb \mem~15 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][112]~q ),
	.datac(!in_data_reg_112),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~15 .extended_lut = "off";
defparam \mem~15 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~15 .shared_arith = "off";

dffeas \mem[1][113] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][113]~q ),
	.prn(vcc));
defparam \mem[1][113] .is_wysiwyg = "true";
defparam \mem[1][113] .power_up = "low";

cyclonev_lcell_comb \mem~16 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][113]~q ),
	.datac(!in_data_reg_113),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~16 .extended_lut = "off";
defparam \mem~16 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~16 .shared_arith = "off";

dffeas \mem[1][114] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][114]~q ),
	.prn(vcc));
defparam \mem[1][114] .is_wysiwyg = "true";
defparam \mem[1][114] .power_up = "low";

cyclonev_lcell_comb \mem~17 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][114]~q ),
	.datac(!in_data_reg_114),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~17 .extended_lut = "off";
defparam \mem~17 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~17 .shared_arith = "off";

dffeas \mem[1][115] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][115]~q ),
	.prn(vcc));
defparam \mem[1][115] .is_wysiwyg = "true";
defparam \mem[1][115] .power_up = "low";

cyclonev_lcell_comb \mem~18 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][115]~q ),
	.datac(!in_data_reg_115),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~18 .extended_lut = "off";
defparam \mem~18 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~18 .shared_arith = "off";

dffeas \mem[1][116] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][116]~q ),
	.prn(vcc));
defparam \mem[1][116] .is_wysiwyg = "true";
defparam \mem[1][116] .power_up = "low";

cyclonev_lcell_comb \mem~19 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][116]~q ),
	.datac(!in_data_reg_116),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~19 .extended_lut = "off";
defparam \mem~19 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~19 .shared_arith = "off";

endmodule

module spw_babasu_altera_avalon_sc_fifo_14 (
	read_latency_shift_reg_0,
	mem_used_0,
	mem_129_0,
	mem_used_01,
	av_readdata_pre_0,
	mem_0_0,
	reset,
	WideOr0,
	clk)/* synthesis synthesis_greybox=0 */;
input 	read_latency_shift_reg_0;
output 	mem_used_0;
input 	mem_129_0;
input 	mem_used_01;
input 	av_readdata_pre_0;
output 	mem_0_0;
input 	reset;
input 	WideOr0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~q ;
wire \mem_used[0]~0_combout ;
wire \mem[1][0]~q ;
wire \mem~0_combout ;
wire \mem[0][0]~1_combout ;


dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][0] (
	.clk(clk),
	.d(\mem[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_0_0),
	.prn(vcc));
defparam \mem[0][0] .is_wysiwyg = "true";
defparam \mem[0][0] .power_up = "low";

cyclonev_lcell_comb \read~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_129_0),
	.datad(!mem_used_01),
	.datae(!WideOr0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h0000777000007770;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!\mem_used[1]~q ),
	.datad(!\read~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'h1F001F001F001F00;
defparam \mem_used[1]~1 .shared_arith = "off";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[1]~q ),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!\mem_used[1]~q ),
	.datad(!\read~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~0 .extended_lut = "off";
defparam \mem_used[0]~0 .lut_mask = 64'h731F731F731F731F;
defparam \mem_used[0]~0 .shared_arith = "off";

dffeas \mem[1][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][0]~q ),
	.prn(vcc));
defparam \mem[1][0] .is_wysiwyg = "true";
defparam \mem[1][0] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!av_readdata_pre_0),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h4747474747474747;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \mem[0][0]~1 (
	.dataa(!mem_used_0),
	.datab(!mem_0_0),
	.datac(!\read~0_combout ),
	.datad(!\mem~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem[0][0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem[0][0]~1 .extended_lut = "off";
defparam \mem[0][0]~1 .lut_mask = 64'h10BF10BF10BF10BF;
defparam \mem[0][0]~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_avalon_sc_fifo_15 (
	out_valid_reg,
	mem_used_1,
	WideOr0,
	in_data_reg_68,
	stateST_UNCOMP_WR_SUBBURST,
	mem_129_0,
	mem_used_0,
	mem_68_0,
	mem_66_0,
	comb,
	mem_130_0,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	mem_105_0,
	mem_106_0,
	mem_107_0,
	mem_108_0,
	mem_109_0,
	mem_110_0,
	mem_111_0,
	mem_112_0,
	mem_113_0,
	mem_114_0,
	mem_115_0,
	mem_116_0,
	reset,
	nxt_out_eop,
	last_packet_beat,
	WideOr01,
	read,
	cp_ready,
	in_data_reg_69,
	rf_source_valid,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_6,
	sink_ready,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	clk)/* synthesis synthesis_greybox=0 */;
input 	out_valid_reg;
output 	mem_used_1;
input 	WideOr0;
input 	in_data_reg_68;
input 	stateST_UNCOMP_WR_SUBBURST;
output 	mem_129_0;
output 	mem_used_0;
output 	mem_68_0;
output 	mem_66_0;
input 	comb;
output 	mem_130_0;
output 	mem_78_0;
output 	mem_77_0;
output 	mem_76_0;
output 	mem_75_0;
output 	mem_74_0;
output 	mem_105_0;
output 	mem_106_0;
output 	mem_107_0;
output 	mem_108_0;
output 	mem_109_0;
output 	mem_110_0;
output 	mem_111_0;
output 	mem_112_0;
output 	mem_113_0;
output 	mem_114_0;
output 	mem_115_0;
output 	mem_116_0;
input 	reset;
input 	nxt_out_eop;
input 	last_packet_beat;
input 	WideOr01;
output 	read;
input 	cp_ready;
input 	in_data_reg_69;
input 	rf_source_valid;
input 	out_byte_cnt_reg_2;
input 	out_uncomp_byte_cnt_reg_4;
input 	out_uncomp_byte_cnt_reg_3;
input 	out_uncomp_byte_cnt_reg_2;
input 	out_uncomp_byte_cnt_reg_5;
input 	out_uncomp_byte_cnt_reg_6;
input 	sink_ready;
input 	in_data_reg_105;
input 	in_data_reg_106;
input 	in_data_reg_107;
input 	in_data_reg_108;
input 	in_data_reg_109;
input 	in_data_reg_110;
input 	in_data_reg_111;
input 	in_data_reg_112;
input 	in_data_reg_113;
input 	in_data_reg_114;
input 	in_data_reg_115;
input 	in_data_reg_116;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \write~0_combout ;
wire \mem_used[1]~0_combout ;
wire \mem[1][129]~q ;
wire \mem~20_combout ;
wire \always0~0_combout ;
wire \mem_used[0]~1_combout ;
wire \mem[1][68]~q ;
wire \mem~0_combout ;
wire \mem[1][66]~q ;
wire \mem~1_combout ;
wire \mem[1][130]~q ;
wire \mem~2_combout ;
wire \mem[1][78]~q ;
wire \mem~3_combout ;
wire \mem[1][77]~q ;
wire \mem~4_combout ;
wire \mem[1][76]~q ;
wire \mem~5_combout ;
wire \mem[1][75]~q ;
wire \mem~6_combout ;
wire \mem[1][74]~q ;
wire \mem~7_combout ;
wire \mem[1][105]~q ;
wire \mem~8_combout ;
wire \mem[1][106]~q ;
wire \mem~9_combout ;
wire \mem[1][107]~q ;
wire \mem~10_combout ;
wire \mem[1][108]~q ;
wire \mem~11_combout ;
wire \mem[1][109]~q ;
wire \mem~12_combout ;
wire \mem[1][110]~q ;
wire \mem~13_combout ;
wire \mem[1][111]~q ;
wire \mem~14_combout ;
wire \mem[1][112]~q ;
wire \mem~15_combout ;
wire \mem[1][113]~q ;
wire \mem~16_combout ;
wire \mem[1][114]~q ;
wire \mem~17_combout ;
wire \mem[1][115]~q ;
wire \mem~18_combout ;
wire \mem[1][116]~q ;
wire \mem~19_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][129] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_129_0),
	.prn(vcc));
defparam \mem[0][129] .is_wysiwyg = "true";
defparam \mem[0][129] .power_up = "low";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][68] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_68_0),
	.prn(vcc));
defparam \mem[0][68] .is_wysiwyg = "true";
defparam \mem[0][68] .power_up = "low";

dffeas \mem[0][66] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_66_0),
	.prn(vcc));
defparam \mem[0][66] .is_wysiwyg = "true";
defparam \mem[0][66] .power_up = "low";

dffeas \mem[0][130] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_130_0),
	.prn(vcc));
defparam \mem[0][130] .is_wysiwyg = "true";
defparam \mem[0][130] .power_up = "low";

dffeas \mem[0][78] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_78_0),
	.prn(vcc));
defparam \mem[0][78] .is_wysiwyg = "true";
defparam \mem[0][78] .power_up = "low";

dffeas \mem[0][77] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_77_0),
	.prn(vcc));
defparam \mem[0][77] .is_wysiwyg = "true";
defparam \mem[0][77] .power_up = "low";

dffeas \mem[0][76] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_76_0),
	.prn(vcc));
defparam \mem[0][76] .is_wysiwyg = "true";
defparam \mem[0][76] .power_up = "low";

dffeas \mem[0][75] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_75_0),
	.prn(vcc));
defparam \mem[0][75] .is_wysiwyg = "true";
defparam \mem[0][75] .power_up = "low";

dffeas \mem[0][74] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_74_0),
	.prn(vcc));
defparam \mem[0][74] .is_wysiwyg = "true";
defparam \mem[0][74] .power_up = "low";

dffeas \mem[0][105] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_105_0),
	.prn(vcc));
defparam \mem[0][105] .is_wysiwyg = "true";
defparam \mem[0][105] .power_up = "low";

dffeas \mem[0][106] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_106_0),
	.prn(vcc));
defparam \mem[0][106] .is_wysiwyg = "true";
defparam \mem[0][106] .power_up = "low";

dffeas \mem[0][107] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_107_0),
	.prn(vcc));
defparam \mem[0][107] .is_wysiwyg = "true";
defparam \mem[0][107] .power_up = "low";

dffeas \mem[0][108] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_108_0),
	.prn(vcc));
defparam \mem[0][108] .is_wysiwyg = "true";
defparam \mem[0][108] .power_up = "low";

dffeas \mem[0][109] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_109_0),
	.prn(vcc));
defparam \mem[0][109] .is_wysiwyg = "true";
defparam \mem[0][109] .power_up = "low";

dffeas \mem[0][110] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_110_0),
	.prn(vcc));
defparam \mem[0][110] .is_wysiwyg = "true";
defparam \mem[0][110] .power_up = "low";

dffeas \mem[0][111] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_111_0),
	.prn(vcc));
defparam \mem[0][111] .is_wysiwyg = "true";
defparam \mem[0][111] .power_up = "low";

dffeas \mem[0][112] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_112_0),
	.prn(vcc));
defparam \mem[0][112] .is_wysiwyg = "true";
defparam \mem[0][112] .power_up = "low";

dffeas \mem[0][113] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_113_0),
	.prn(vcc));
defparam \mem[0][113] .is_wysiwyg = "true";
defparam \mem[0][113] .power_up = "low";

dffeas \mem[0][114] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_114_0),
	.prn(vcc));
defparam \mem[0][114] .is_wysiwyg = "true";
defparam \mem[0][114] .power_up = "low";

dffeas \mem[0][115] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_115_0),
	.prn(vcc));
defparam \mem[0][115] .is_wysiwyg = "true";
defparam \mem[0][115] .power_up = "low";

dffeas \mem[0][116] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_116_0),
	.prn(vcc));
defparam \mem[0][116] .is_wysiwyg = "true";
defparam \mem[0][116] .power_up = "low";

cyclonev_lcell_comb \read~0 (
	.dataa(!comb),
	.datab(!WideOr01),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h1111111111111111;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \write~0 (
	.dataa(!mem_used_1),
	.datab(!WideOr0),
	.datac(!cp_ready),
	.datad(!rf_source_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'h008A008A008A008A;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!last_packet_beat),
	.datad(!read),
	.datae(!\write~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'h5505335355053353;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][129] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][129]~q ),
	.prn(vcc));
defparam \mem[1][129] .is_wysiwyg = "true";
defparam \mem[1][129] .power_up = "low";

cyclonev_lcell_comb \mem~20 (
	.dataa(!WideOr0),
	.datab(!out_valid_reg),
	.datac(!\mem[1][129]~q ),
	.datad(!in_data_reg_68),
	.datae(!mem_used_1),
	.dataf(!nxt_out_eop),
	.datag(!in_data_reg_69),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~20 .extended_lut = "on";
defparam \mem~20 .lut_mask = 64'h02020F0F02330F0F;
defparam \mem~20 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!mem_used_0),
	.datab(!sink_ready),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!\write~0_combout ),
	.datad(!sink_ready),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'h3F1F3F1F3F1F3F1F;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem[1][68] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][68]~q ),
	.prn(vcc));
defparam \mem[1][68] .is_wysiwyg = "true";
defparam \mem[1][68] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!mem_used_1),
	.datab(!in_data_reg_68),
	.datac(!\mem[1][68]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h2727272727272727;
defparam \mem~0 .shared_arith = "off";

dffeas \mem[1][66] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][66]~q ),
	.prn(vcc));
defparam \mem[1][66] .is_wysiwyg = "true";
defparam \mem[1][66] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!mem_used_1),
	.datab(!in_data_reg_69),
	.datac(!\mem[1][66]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h2727272727272727;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[1][130] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][130]~q ),
	.prn(vcc));
defparam \mem[1][130] .is_wysiwyg = "true";
defparam \mem[1][130] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!mem_used_1),
	.datab(!nxt_out_eop),
	.datac(!\mem[1][130]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h2727272727272727;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[1][78] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][78]~q ),
	.prn(vcc));
defparam \mem[1][78] .is_wysiwyg = "true";
defparam \mem[1][78] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_6),
	.datad(!\mem[1][78]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h0257025702570257;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][77] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][77]~q ),
	.prn(vcc));
defparam \mem[1][77] .is_wysiwyg = "true";
defparam \mem[1][77] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\mem[1][77]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h0257025702570257;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][76] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][76]~q ),
	.prn(vcc));
defparam \mem[1][76] .is_wysiwyg = "true";
defparam \mem[1][76] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!\mem[1][76]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h0257025702570257;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][75] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][75]~q ),
	.prn(vcc));
defparam \mem[1][75] .is_wysiwyg = "true";
defparam \mem[1][75] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\mem[1][75]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h0257025702570257;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[1][74] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][74]~q ),
	.prn(vcc));
defparam \mem[1][74] .is_wysiwyg = "true";
defparam \mem[1][74] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_byte_cnt_reg_2),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(!\mem[1][74]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h082A5D7F082A5D7F;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[1][105] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][105]~q ),
	.prn(vcc));
defparam \mem[1][105] .is_wysiwyg = "true";
defparam \mem[1][105] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][105]~q ),
	.datac(!in_data_reg_105),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~8 .shared_arith = "off";

dffeas \mem[1][106] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][106]~q ),
	.prn(vcc));
defparam \mem[1][106] .is_wysiwyg = "true";
defparam \mem[1][106] .power_up = "low";

cyclonev_lcell_comb \mem~9 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][106]~q ),
	.datac(!in_data_reg_106),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~9 .extended_lut = "off";
defparam \mem~9 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~9 .shared_arith = "off";

dffeas \mem[1][107] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][107]~q ),
	.prn(vcc));
defparam \mem[1][107] .is_wysiwyg = "true";
defparam \mem[1][107] .power_up = "low";

cyclonev_lcell_comb \mem~10 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][107]~q ),
	.datac(!in_data_reg_107),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~10 .extended_lut = "off";
defparam \mem~10 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~10 .shared_arith = "off";

dffeas \mem[1][108] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][108]~q ),
	.prn(vcc));
defparam \mem[1][108] .is_wysiwyg = "true";
defparam \mem[1][108] .power_up = "low";

cyclonev_lcell_comb \mem~11 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][108]~q ),
	.datac(!in_data_reg_108),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~11 .extended_lut = "off";
defparam \mem~11 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~11 .shared_arith = "off";

dffeas \mem[1][109] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][109]~q ),
	.prn(vcc));
defparam \mem[1][109] .is_wysiwyg = "true";
defparam \mem[1][109] .power_up = "low";

cyclonev_lcell_comb \mem~12 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][109]~q ),
	.datac(!in_data_reg_109),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~12 .extended_lut = "off";
defparam \mem~12 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~12 .shared_arith = "off";

dffeas \mem[1][110] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][110]~q ),
	.prn(vcc));
defparam \mem[1][110] .is_wysiwyg = "true";
defparam \mem[1][110] .power_up = "low";

cyclonev_lcell_comb \mem~13 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][110]~q ),
	.datac(!in_data_reg_110),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~13 .extended_lut = "off";
defparam \mem~13 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~13 .shared_arith = "off";

dffeas \mem[1][111] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][111]~q ),
	.prn(vcc));
defparam \mem[1][111] .is_wysiwyg = "true";
defparam \mem[1][111] .power_up = "low";

cyclonev_lcell_comb \mem~14 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][111]~q ),
	.datac(!in_data_reg_111),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~14 .extended_lut = "off";
defparam \mem~14 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~14 .shared_arith = "off";

dffeas \mem[1][112] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][112]~q ),
	.prn(vcc));
defparam \mem[1][112] .is_wysiwyg = "true";
defparam \mem[1][112] .power_up = "low";

cyclonev_lcell_comb \mem~15 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][112]~q ),
	.datac(!in_data_reg_112),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~15 .extended_lut = "off";
defparam \mem~15 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~15 .shared_arith = "off";

dffeas \mem[1][113] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][113]~q ),
	.prn(vcc));
defparam \mem[1][113] .is_wysiwyg = "true";
defparam \mem[1][113] .power_up = "low";

cyclonev_lcell_comb \mem~16 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][113]~q ),
	.datac(!in_data_reg_113),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~16 .extended_lut = "off";
defparam \mem~16 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~16 .shared_arith = "off";

dffeas \mem[1][114] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][114]~q ),
	.prn(vcc));
defparam \mem[1][114] .is_wysiwyg = "true";
defparam \mem[1][114] .power_up = "low";

cyclonev_lcell_comb \mem~17 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][114]~q ),
	.datac(!in_data_reg_114),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~17 .extended_lut = "off";
defparam \mem~17 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~17 .shared_arith = "off";

dffeas \mem[1][115] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][115]~q ),
	.prn(vcc));
defparam \mem[1][115] .is_wysiwyg = "true";
defparam \mem[1][115] .power_up = "low";

cyclonev_lcell_comb \mem~18 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][115]~q ),
	.datac(!in_data_reg_115),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~18 .extended_lut = "off";
defparam \mem~18 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~18 .shared_arith = "off";

dffeas \mem[1][116] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][116]~q ),
	.prn(vcc));
defparam \mem[1][116] .is_wysiwyg = "true";
defparam \mem[1][116] .power_up = "low";

cyclonev_lcell_comb \mem~19 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][116]~q ),
	.datac(!in_data_reg_116),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~19 .extended_lut = "off";
defparam \mem~19 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~19 .shared_arith = "off";

endmodule

module spw_babasu_altera_avalon_sc_fifo_16 (
	h2f_RREADY_0,
	read_latency_shift_reg_0,
	mem_used_0,
	empty1,
	av_readdata_pre_0,
	mem_0_0,
	reset,
	clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_RREADY_0;
input 	read_latency_shift_reg_0;
output 	mem_used_0;
output 	empty1;
input 	av_readdata_pre_0;
output 	mem_0_0;
input 	reset;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[1]~1_combout ;
wire \mem_used[1]~q ;
wire \mem_used[0]~0_combout ;
wire \mem[1][0]~q ;
wire \mem~0_combout ;
wire \mem[0][0]~1_combout ;


dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb empty(
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(empty1),
	.sumout(),
	.cout(),
	.shareout());
defparam empty.extended_lut = "off";
defparam empty.lut_mask = 64'h8888888888888888;
defparam empty.shared_arith = "off";

dffeas \mem[0][0] (
	.clk(clk),
	.d(\mem[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_0_0),
	.prn(vcc));
defparam \mem[0][0] .is_wysiwyg = "true";
defparam \mem[0][0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!h2f_RREADY_0),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem_used[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'h02EA02EA02EA02EA;
defparam \mem_used[1]~1 .shared_arith = "off";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[1]~q ),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~0 (
	.dataa(!h2f_RREADY_0),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem_used[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~0 .extended_lut = "off";
defparam \mem_used[0]~0 .lut_mask = 64'h2B1F2B1F2B1F2B1F;
defparam \mem_used[0]~0 .shared_arith = "off";

dffeas \mem[1][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][0]~q ),
	.prn(vcc));
defparam \mem[1][0] .is_wysiwyg = "true";
defparam \mem[1][0] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!av_readdata_pre_0),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h4747474747474747;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \mem[0][0]~1 (
	.dataa(!h2f_RREADY_0),
	.datab(!mem_used_0),
	.datac(!mem_0_0),
	.datad(!\mem~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem[0][0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem[0][0]~1 .extended_lut = "off";
defparam \mem[0][0]~1 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \mem[0][0]~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_avalon_sc_fifo_17 (
	h2f_RREADY_0,
	waitrequest_reset_override,
	mem_used_1,
	in_data_reg_69,
	wait_latency_counter_1,
	wait_latency_counter_0,
	nxt_out_eop,
	out_valid_reg,
	stateST_UNCOMP_WR_SUBBURST,
	mem_130_0,
	empty,
	mem_66_0,
	mem_used_0,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	mem_105_0,
	mem_106_0,
	mem_107_0,
	mem_108_0,
	mem_109_0,
	mem_110_0,
	mem_111_0,
	mem_112_0,
	mem_113_0,
	mem_114_0,
	mem_115_0,
	mem_116_0,
	reset,
	last_packet_beat,
	write,
	write1,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_6,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_RREADY_0;
input 	waitrequest_reset_override;
output 	mem_used_1;
input 	in_data_reg_69;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	nxt_out_eop;
input 	out_valid_reg;
input 	stateST_UNCOMP_WR_SUBBURST;
output 	mem_130_0;
input 	empty;
output 	mem_66_0;
output 	mem_used_0;
output 	mem_78_0;
output 	mem_77_0;
output 	mem_76_0;
output 	mem_75_0;
output 	mem_74_0;
output 	mem_105_0;
output 	mem_106_0;
output 	mem_107_0;
output 	mem_108_0;
output 	mem_109_0;
output 	mem_110_0;
output 	mem_111_0;
output 	mem_112_0;
output 	mem_113_0;
output 	mem_114_0;
output 	mem_115_0;
output 	mem_116_0;
input 	reset;
input 	last_packet_beat;
output 	write;
output 	write1;
input 	out_byte_cnt_reg_2;
input 	out_uncomp_byte_cnt_reg_5;
input 	out_uncomp_byte_cnt_reg_4;
input 	out_uncomp_byte_cnt_reg_3;
input 	out_uncomp_byte_cnt_reg_2;
input 	out_uncomp_byte_cnt_reg_6;
input 	in_data_reg_105;
input 	in_data_reg_106;
input 	in_data_reg_107;
input 	in_data_reg_108;
input 	in_data_reg_109;
input 	in_data_reg_110;
input 	in_data_reg_111;
input 	in_data_reg_112;
input 	in_data_reg_113;
input 	in_data_reg_114;
input 	in_data_reg_115;
input 	in_data_reg_116;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read~0_combout ;
wire \mem_used[1]~0_combout ;
wire \mem[1][130]~q ;
wire \mem~0_combout ;
wire \always0~0_combout ;
wire \mem[1][69]~q ;
wire \mem~1_combout ;
wire \mem_used[0]~1_combout ;
wire \mem[1][78]~q ;
wire \mem~2_combout ;
wire \mem[1][77]~q ;
wire \mem~3_combout ;
wire \mem[1][76]~q ;
wire \mem~4_combout ;
wire \mem[1][75]~q ;
wire \mem~5_combout ;
wire \mem[1][74]~q ;
wire \mem~6_combout ;
wire \mem[1][105]~q ;
wire \mem~7_combout ;
wire \mem[1][106]~q ;
wire \mem~8_combout ;
wire \mem[1][107]~q ;
wire \mem~9_combout ;
wire \mem[1][108]~q ;
wire \mem~10_combout ;
wire \mem[1][109]~q ;
wire \mem~11_combout ;
wire \mem[1][110]~q ;
wire \mem~12_combout ;
wire \mem[1][111]~q ;
wire \mem~13_combout ;
wire \mem[1][112]~q ;
wire \mem~14_combout ;
wire \mem[1][113]~q ;
wire \mem~15_combout ;
wire \mem[1][114]~q ;
wire \mem~16_combout ;
wire \mem[1][115]~q ;
wire \mem~17_combout ;
wire \mem[1][116]~q ;
wire \mem~18_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][130] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_130_0),
	.prn(vcc));
defparam \mem[0][130] .is_wysiwyg = "true";
defparam \mem[0][130] .power_up = "low";

dffeas \mem[0][66] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_66_0),
	.prn(vcc));
defparam \mem[0][66] .is_wysiwyg = "true";
defparam \mem[0][66] .power_up = "low";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][78] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_78_0),
	.prn(vcc));
defparam \mem[0][78] .is_wysiwyg = "true";
defparam \mem[0][78] .power_up = "low";

dffeas \mem[0][77] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_77_0),
	.prn(vcc));
defparam \mem[0][77] .is_wysiwyg = "true";
defparam \mem[0][77] .power_up = "low";

dffeas \mem[0][76] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_76_0),
	.prn(vcc));
defparam \mem[0][76] .is_wysiwyg = "true";
defparam \mem[0][76] .power_up = "low";

dffeas \mem[0][75] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_75_0),
	.prn(vcc));
defparam \mem[0][75] .is_wysiwyg = "true";
defparam \mem[0][75] .power_up = "low";

dffeas \mem[0][74] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_74_0),
	.prn(vcc));
defparam \mem[0][74] .is_wysiwyg = "true";
defparam \mem[0][74] .power_up = "low";

dffeas \mem[0][105] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_105_0),
	.prn(vcc));
defparam \mem[0][105] .is_wysiwyg = "true";
defparam \mem[0][105] .power_up = "low";

dffeas \mem[0][106] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_106_0),
	.prn(vcc));
defparam \mem[0][106] .is_wysiwyg = "true";
defparam \mem[0][106] .power_up = "low";

dffeas \mem[0][107] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_107_0),
	.prn(vcc));
defparam \mem[0][107] .is_wysiwyg = "true";
defparam \mem[0][107] .power_up = "low";

dffeas \mem[0][108] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_108_0),
	.prn(vcc));
defparam \mem[0][108] .is_wysiwyg = "true";
defparam \mem[0][108] .power_up = "low";

dffeas \mem[0][109] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_109_0),
	.prn(vcc));
defparam \mem[0][109] .is_wysiwyg = "true";
defparam \mem[0][109] .power_up = "low";

dffeas \mem[0][110] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_110_0),
	.prn(vcc));
defparam \mem[0][110] .is_wysiwyg = "true";
defparam \mem[0][110] .power_up = "low";

dffeas \mem[0][111] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_111_0),
	.prn(vcc));
defparam \mem[0][111] .is_wysiwyg = "true";
defparam \mem[0][111] .power_up = "low";

dffeas \mem[0][112] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_112_0),
	.prn(vcc));
defparam \mem[0][112] .is_wysiwyg = "true";
defparam \mem[0][112] .power_up = "low";

dffeas \mem[0][113] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_113_0),
	.prn(vcc));
defparam \mem[0][113] .is_wysiwyg = "true";
defparam \mem[0][113] .power_up = "low";

dffeas \mem[0][114] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_114_0),
	.prn(vcc));
defparam \mem[0][114] .is_wysiwyg = "true";
defparam \mem[0][114] .power_up = "low";

dffeas \mem[0][115] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_115_0),
	.prn(vcc));
defparam \mem[0][115] .is_wysiwyg = "true";
defparam \mem[0][115] .power_up = "low";

dffeas \mem[0][116] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_116_0),
	.prn(vcc));
defparam \mem[0][116] .is_wysiwyg = "true";
defparam \mem[0][116] .power_up = "low";

cyclonev_lcell_comb \write~0 (
	.dataa(!waitrequest_reset_override),
	.datab(!in_data_reg_69),
	.datac(!mem_used_1),
	.datad(!out_valid_reg),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'h0010001000100010;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \write~1 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!write),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write1),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~1 .extended_lut = "off";
defparam \write~1 .lut_mask = 64'h0202020202020202;
defparam \write~1 .shared_arith = "off";

cyclonev_lcell_comb \read~0 (
	.dataa(!h2f_RREADY_0),
	.datab(!empty),
	.datac(!last_packet_beat),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h4040404040404040;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!\read~0_combout ),
	.datad(!write1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'h5431543154315431;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][130] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][130]~q ),
	.prn(vcc));
defparam \mem[1][130] .is_wysiwyg = "true";
defparam \mem[1][130] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!mem_used_1),
	.datab(!nxt_out_eop),
	.datac(!\mem[1][130]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h2727272727272727;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!mem_used_0),
	.datab(!\read~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \always0~0 .shared_arith = "off";

dffeas \mem[1][69] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][69]~q ),
	.prn(vcc));
defparam \mem[1][69] .is_wysiwyg = "true";
defparam \mem[1][69] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!in_data_reg_69),
	.datab(!mem_used_1),
	.datac(!\mem[1][69]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h4747474747474747;
defparam \mem~1 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!\read~0_combout ),
	.datad(!write1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'h31FF31FF31FF31FF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem[1][78] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][78]~q ),
	.prn(vcc));
defparam \mem[1][78] .is_wysiwyg = "true";
defparam \mem[1][78] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_6),
	.datad(!\mem[1][78]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h0257025702570257;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[1][77] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][77]~q ),
	.prn(vcc));
defparam \mem[1][77] .is_wysiwyg = "true";
defparam \mem[1][77] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\mem[1][77]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h0257025702570257;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][76] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][76]~q ),
	.prn(vcc));
defparam \mem[1][76] .is_wysiwyg = "true";
defparam \mem[1][76] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!\mem[1][76]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h0257025702570257;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][75] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][75]~q ),
	.prn(vcc));
defparam \mem[1][75] .is_wysiwyg = "true";
defparam \mem[1][75] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\mem[1][75]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h0257025702570257;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][74] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][74]~q ),
	.prn(vcc));
defparam \mem[1][74] .is_wysiwyg = "true";
defparam \mem[1][74] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_byte_cnt_reg_2),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(!\mem[1][74]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h082A5D7F082A5D7F;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[1][105] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][105]~q ),
	.prn(vcc));
defparam \mem[1][105] .is_wysiwyg = "true";
defparam \mem[1][105] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][105]~q ),
	.datac(!in_data_reg_105),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[1][106] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][106]~q ),
	.prn(vcc));
defparam \mem[1][106] .is_wysiwyg = "true";
defparam \mem[1][106] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][106]~q ),
	.datac(!in_data_reg_106),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~8 .shared_arith = "off";

dffeas \mem[1][107] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][107]~q ),
	.prn(vcc));
defparam \mem[1][107] .is_wysiwyg = "true";
defparam \mem[1][107] .power_up = "low";

cyclonev_lcell_comb \mem~9 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][107]~q ),
	.datac(!in_data_reg_107),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~9 .extended_lut = "off";
defparam \mem~9 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~9 .shared_arith = "off";

dffeas \mem[1][108] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][108]~q ),
	.prn(vcc));
defparam \mem[1][108] .is_wysiwyg = "true";
defparam \mem[1][108] .power_up = "low";

cyclonev_lcell_comb \mem~10 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][108]~q ),
	.datac(!in_data_reg_108),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~10 .extended_lut = "off";
defparam \mem~10 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~10 .shared_arith = "off";

dffeas \mem[1][109] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][109]~q ),
	.prn(vcc));
defparam \mem[1][109] .is_wysiwyg = "true";
defparam \mem[1][109] .power_up = "low";

cyclonev_lcell_comb \mem~11 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][109]~q ),
	.datac(!in_data_reg_109),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~11 .extended_lut = "off";
defparam \mem~11 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~11 .shared_arith = "off";

dffeas \mem[1][110] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][110]~q ),
	.prn(vcc));
defparam \mem[1][110] .is_wysiwyg = "true";
defparam \mem[1][110] .power_up = "low";

cyclonev_lcell_comb \mem~12 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][110]~q ),
	.datac(!in_data_reg_110),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~12 .extended_lut = "off";
defparam \mem~12 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~12 .shared_arith = "off";

dffeas \mem[1][111] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][111]~q ),
	.prn(vcc));
defparam \mem[1][111] .is_wysiwyg = "true";
defparam \mem[1][111] .power_up = "low";

cyclonev_lcell_comb \mem~13 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][111]~q ),
	.datac(!in_data_reg_111),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~13 .extended_lut = "off";
defparam \mem~13 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~13 .shared_arith = "off";

dffeas \mem[1][112] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][112]~q ),
	.prn(vcc));
defparam \mem[1][112] .is_wysiwyg = "true";
defparam \mem[1][112] .power_up = "low";

cyclonev_lcell_comb \mem~14 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][112]~q ),
	.datac(!in_data_reg_112),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~14 .extended_lut = "off";
defparam \mem~14 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~14 .shared_arith = "off";

dffeas \mem[1][113] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][113]~q ),
	.prn(vcc));
defparam \mem[1][113] .is_wysiwyg = "true";
defparam \mem[1][113] .power_up = "low";

cyclonev_lcell_comb \mem~15 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][113]~q ),
	.datac(!in_data_reg_113),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~15 .extended_lut = "off";
defparam \mem~15 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~15 .shared_arith = "off";

dffeas \mem[1][114] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][114]~q ),
	.prn(vcc));
defparam \mem[1][114] .is_wysiwyg = "true";
defparam \mem[1][114] .power_up = "low";

cyclonev_lcell_comb \mem~16 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][114]~q ),
	.datac(!in_data_reg_114),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~16 .extended_lut = "off";
defparam \mem~16 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~16 .shared_arith = "off";

dffeas \mem[1][115] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][115]~q ),
	.prn(vcc));
defparam \mem[1][115] .is_wysiwyg = "true";
defparam \mem[1][115] .power_up = "low";

cyclonev_lcell_comb \mem~17 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][115]~q ),
	.datac(!in_data_reg_115),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~17 .extended_lut = "off";
defparam \mem~17 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~17 .shared_arith = "off";

dffeas \mem[1][116] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][116]~q ),
	.prn(vcc));
defparam \mem[1][116] .is_wysiwyg = "true";
defparam \mem[1][116] .power_up = "low";

cyclonev_lcell_comb \mem~18 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][116]~q ),
	.datac(!in_data_reg_116),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~18 .extended_lut = "off";
defparam \mem~18 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~18 .shared_arith = "off";

endmodule

module spw_babasu_altera_avalon_sc_fifo_18 (
	read_latency_shift_reg_0,
	mem_used_0,
	mem_129_0,
	mem_used_01,
	av_readdata_pre_0,
	mem_0_0,
	reset,
	WideOr0,
	clk)/* synthesis synthesis_greybox=0 */;
input 	read_latency_shift_reg_0;
output 	mem_used_0;
input 	mem_129_0;
input 	mem_used_01;
input 	av_readdata_pre_0;
output 	mem_0_0;
input 	reset;
input 	WideOr0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~q ;
wire \mem_used[0]~0_combout ;
wire \mem[1][0]~q ;
wire \mem~0_combout ;
wire \mem[0][0]~1_combout ;


dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][0] (
	.clk(clk),
	.d(\mem[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_0_0),
	.prn(vcc));
defparam \mem[0][0] .is_wysiwyg = "true";
defparam \mem[0][0] .power_up = "low";

cyclonev_lcell_comb \read~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_129_0),
	.datad(!mem_used_01),
	.datae(!WideOr0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h0000777000007770;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!\mem_used[1]~q ),
	.datad(!\read~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'h1F001F001F001F00;
defparam \mem_used[1]~1 .shared_arith = "off";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[1]~q ),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!\mem_used[1]~q ),
	.datad(!\read~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~0 .extended_lut = "off";
defparam \mem_used[0]~0 .lut_mask = 64'h731F731F731F731F;
defparam \mem_used[0]~0 .shared_arith = "off";

dffeas \mem[1][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][0]~q ),
	.prn(vcc));
defparam \mem[1][0] .is_wysiwyg = "true";
defparam \mem[1][0] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!av_readdata_pre_0),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h4747474747474747;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \mem[0][0]~1 (
	.dataa(!mem_used_0),
	.datab(!mem_0_0),
	.datac(!\read~0_combout ),
	.datad(!\mem~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem[0][0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem[0][0]~1 .extended_lut = "off";
defparam \mem[0][0]~1 .lut_mask = 64'h10BF10BF10BF10BF;
defparam \mem[0][0]~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_avalon_sc_fifo_19 (
	out_valid_reg,
	mem_used_1,
	WideOr0,
	in_data_reg_68,
	stateST_UNCOMP_WR_SUBBURST,
	mem_129_0,
	mem_used_0,
	mem_68_0,
	mem_66_0,
	comb,
	mem_130_0,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	mem_105_0,
	mem_106_0,
	mem_107_0,
	mem_108_0,
	mem_109_0,
	mem_110_0,
	mem_111_0,
	mem_112_0,
	mem_113_0,
	mem_114_0,
	mem_115_0,
	mem_116_0,
	reset,
	nxt_out_eop,
	last_packet_beat,
	WideOr01,
	read,
	cp_ready,
	in_data_reg_69,
	rf_source_valid,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_6,
	sink_ready,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	clk)/* synthesis synthesis_greybox=0 */;
input 	out_valid_reg;
output 	mem_used_1;
input 	WideOr0;
input 	in_data_reg_68;
input 	stateST_UNCOMP_WR_SUBBURST;
output 	mem_129_0;
output 	mem_used_0;
output 	mem_68_0;
output 	mem_66_0;
input 	comb;
output 	mem_130_0;
output 	mem_78_0;
output 	mem_77_0;
output 	mem_76_0;
output 	mem_75_0;
output 	mem_74_0;
output 	mem_105_0;
output 	mem_106_0;
output 	mem_107_0;
output 	mem_108_0;
output 	mem_109_0;
output 	mem_110_0;
output 	mem_111_0;
output 	mem_112_0;
output 	mem_113_0;
output 	mem_114_0;
output 	mem_115_0;
output 	mem_116_0;
input 	reset;
input 	nxt_out_eop;
input 	last_packet_beat;
input 	WideOr01;
output 	read;
input 	cp_ready;
input 	in_data_reg_69;
input 	rf_source_valid;
input 	out_byte_cnt_reg_2;
input 	out_uncomp_byte_cnt_reg_5;
input 	out_uncomp_byte_cnt_reg_4;
input 	out_uncomp_byte_cnt_reg_3;
input 	out_uncomp_byte_cnt_reg_2;
input 	out_uncomp_byte_cnt_reg_6;
input 	sink_ready;
input 	in_data_reg_105;
input 	in_data_reg_106;
input 	in_data_reg_107;
input 	in_data_reg_108;
input 	in_data_reg_109;
input 	in_data_reg_110;
input 	in_data_reg_111;
input 	in_data_reg_112;
input 	in_data_reg_113;
input 	in_data_reg_114;
input 	in_data_reg_115;
input 	in_data_reg_116;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \write~0_combout ;
wire \mem_used[1]~0_combout ;
wire \mem[1][129]~q ;
wire \mem~20_combout ;
wire \always0~0_combout ;
wire \mem_used[0]~1_combout ;
wire \mem[1][68]~q ;
wire \mem~0_combout ;
wire \mem[1][69]~q ;
wire \mem~1_combout ;
wire \mem[1][130]~q ;
wire \mem~2_combout ;
wire \mem[1][78]~q ;
wire \mem~3_combout ;
wire \mem[1][77]~q ;
wire \mem~4_combout ;
wire \mem[1][76]~q ;
wire \mem~5_combout ;
wire \mem[1][75]~q ;
wire \mem~6_combout ;
wire \mem[1][74]~q ;
wire \mem~7_combout ;
wire \mem[1][105]~q ;
wire \mem~8_combout ;
wire \mem[1][106]~q ;
wire \mem~9_combout ;
wire \mem[1][107]~q ;
wire \mem~10_combout ;
wire \mem[1][108]~q ;
wire \mem~11_combout ;
wire \mem[1][109]~q ;
wire \mem~12_combout ;
wire \mem[1][110]~q ;
wire \mem~13_combout ;
wire \mem[1][111]~q ;
wire \mem~14_combout ;
wire \mem[1][112]~q ;
wire \mem~15_combout ;
wire \mem[1][113]~q ;
wire \mem~16_combout ;
wire \mem[1][114]~q ;
wire \mem~17_combout ;
wire \mem[1][115]~q ;
wire \mem~18_combout ;
wire \mem[1][116]~q ;
wire \mem~19_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][129] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_129_0),
	.prn(vcc));
defparam \mem[0][129] .is_wysiwyg = "true";
defparam \mem[0][129] .power_up = "low";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][68] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_68_0),
	.prn(vcc));
defparam \mem[0][68] .is_wysiwyg = "true";
defparam \mem[0][68] .power_up = "low";

dffeas \mem[0][66] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_66_0),
	.prn(vcc));
defparam \mem[0][66] .is_wysiwyg = "true";
defparam \mem[0][66] .power_up = "low";

dffeas \mem[0][130] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_130_0),
	.prn(vcc));
defparam \mem[0][130] .is_wysiwyg = "true";
defparam \mem[0][130] .power_up = "low";

dffeas \mem[0][78] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_78_0),
	.prn(vcc));
defparam \mem[0][78] .is_wysiwyg = "true";
defparam \mem[0][78] .power_up = "low";

dffeas \mem[0][77] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_77_0),
	.prn(vcc));
defparam \mem[0][77] .is_wysiwyg = "true";
defparam \mem[0][77] .power_up = "low";

dffeas \mem[0][76] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_76_0),
	.prn(vcc));
defparam \mem[0][76] .is_wysiwyg = "true";
defparam \mem[0][76] .power_up = "low";

dffeas \mem[0][75] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_75_0),
	.prn(vcc));
defparam \mem[0][75] .is_wysiwyg = "true";
defparam \mem[0][75] .power_up = "low";

dffeas \mem[0][74] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_74_0),
	.prn(vcc));
defparam \mem[0][74] .is_wysiwyg = "true";
defparam \mem[0][74] .power_up = "low";

dffeas \mem[0][105] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_105_0),
	.prn(vcc));
defparam \mem[0][105] .is_wysiwyg = "true";
defparam \mem[0][105] .power_up = "low";

dffeas \mem[0][106] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_106_0),
	.prn(vcc));
defparam \mem[0][106] .is_wysiwyg = "true";
defparam \mem[0][106] .power_up = "low";

dffeas \mem[0][107] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_107_0),
	.prn(vcc));
defparam \mem[0][107] .is_wysiwyg = "true";
defparam \mem[0][107] .power_up = "low";

dffeas \mem[0][108] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_108_0),
	.prn(vcc));
defparam \mem[0][108] .is_wysiwyg = "true";
defparam \mem[0][108] .power_up = "low";

dffeas \mem[0][109] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_109_0),
	.prn(vcc));
defparam \mem[0][109] .is_wysiwyg = "true";
defparam \mem[0][109] .power_up = "low";

dffeas \mem[0][110] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_110_0),
	.prn(vcc));
defparam \mem[0][110] .is_wysiwyg = "true";
defparam \mem[0][110] .power_up = "low";

dffeas \mem[0][111] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_111_0),
	.prn(vcc));
defparam \mem[0][111] .is_wysiwyg = "true";
defparam \mem[0][111] .power_up = "low";

dffeas \mem[0][112] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_112_0),
	.prn(vcc));
defparam \mem[0][112] .is_wysiwyg = "true";
defparam \mem[0][112] .power_up = "low";

dffeas \mem[0][113] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_113_0),
	.prn(vcc));
defparam \mem[0][113] .is_wysiwyg = "true";
defparam \mem[0][113] .power_up = "low";

dffeas \mem[0][114] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_114_0),
	.prn(vcc));
defparam \mem[0][114] .is_wysiwyg = "true";
defparam \mem[0][114] .power_up = "low";

dffeas \mem[0][115] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_115_0),
	.prn(vcc));
defparam \mem[0][115] .is_wysiwyg = "true";
defparam \mem[0][115] .power_up = "low";

dffeas \mem[0][116] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_116_0),
	.prn(vcc));
defparam \mem[0][116] .is_wysiwyg = "true";
defparam \mem[0][116] .power_up = "low";

cyclonev_lcell_comb \read~0 (
	.dataa(!comb),
	.datab(!WideOr01),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h1111111111111111;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \write~0 (
	.dataa(!mem_used_1),
	.datab(!WideOr0),
	.datac(!cp_ready),
	.datad(!rf_source_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'h008A008A008A008A;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!last_packet_beat),
	.datad(!read),
	.datae(!\write~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'h5505335355053353;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][129] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][129]~q ),
	.prn(vcc));
defparam \mem[1][129] .is_wysiwyg = "true";
defparam \mem[1][129] .power_up = "low";

cyclonev_lcell_comb \mem~20 (
	.dataa(!WideOr0),
	.datab(!out_valid_reg),
	.datac(!\mem[1][129]~q ),
	.datad(!in_data_reg_68),
	.datae(!mem_used_1),
	.dataf(!nxt_out_eop),
	.datag(!in_data_reg_69),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~20 .extended_lut = "on";
defparam \mem~20 .lut_mask = 64'h02020F0F02330F0F;
defparam \mem~20 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!mem_used_0),
	.datab(!sink_ready),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!\write~0_combout ),
	.datad(!sink_ready),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'h3F1F3F1F3F1F3F1F;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem[1][68] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][68]~q ),
	.prn(vcc));
defparam \mem[1][68] .is_wysiwyg = "true";
defparam \mem[1][68] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!mem_used_1),
	.datab(!in_data_reg_68),
	.datac(!\mem[1][68]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h2727272727272727;
defparam \mem~0 .shared_arith = "off";

dffeas \mem[1][69] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][69]~q ),
	.prn(vcc));
defparam \mem[1][69] .is_wysiwyg = "true";
defparam \mem[1][69] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!mem_used_1),
	.datab(!in_data_reg_69),
	.datac(!\mem[1][69]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h2727272727272727;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[1][130] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][130]~q ),
	.prn(vcc));
defparam \mem[1][130] .is_wysiwyg = "true";
defparam \mem[1][130] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!mem_used_1),
	.datab(!nxt_out_eop),
	.datac(!\mem[1][130]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h2727272727272727;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[1][78] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][78]~q ),
	.prn(vcc));
defparam \mem[1][78] .is_wysiwyg = "true";
defparam \mem[1][78] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_6),
	.datad(!\mem[1][78]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h0257025702570257;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][77] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][77]~q ),
	.prn(vcc));
defparam \mem[1][77] .is_wysiwyg = "true";
defparam \mem[1][77] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\mem[1][77]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h0257025702570257;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][76] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][76]~q ),
	.prn(vcc));
defparam \mem[1][76] .is_wysiwyg = "true";
defparam \mem[1][76] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!\mem[1][76]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h0257025702570257;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][75] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][75]~q ),
	.prn(vcc));
defparam \mem[1][75] .is_wysiwyg = "true";
defparam \mem[1][75] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\mem[1][75]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h0257025702570257;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[1][74] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][74]~q ),
	.prn(vcc));
defparam \mem[1][74] .is_wysiwyg = "true";
defparam \mem[1][74] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_byte_cnt_reg_2),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(!\mem[1][74]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h082A5D7F082A5D7F;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[1][105] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][105]~q ),
	.prn(vcc));
defparam \mem[1][105] .is_wysiwyg = "true";
defparam \mem[1][105] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][105]~q ),
	.datac(!in_data_reg_105),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~8 .shared_arith = "off";

dffeas \mem[1][106] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][106]~q ),
	.prn(vcc));
defparam \mem[1][106] .is_wysiwyg = "true";
defparam \mem[1][106] .power_up = "low";

cyclonev_lcell_comb \mem~9 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][106]~q ),
	.datac(!in_data_reg_106),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~9 .extended_lut = "off";
defparam \mem~9 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~9 .shared_arith = "off";

dffeas \mem[1][107] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][107]~q ),
	.prn(vcc));
defparam \mem[1][107] .is_wysiwyg = "true";
defparam \mem[1][107] .power_up = "low";

cyclonev_lcell_comb \mem~10 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][107]~q ),
	.datac(!in_data_reg_107),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~10 .extended_lut = "off";
defparam \mem~10 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~10 .shared_arith = "off";

dffeas \mem[1][108] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][108]~q ),
	.prn(vcc));
defparam \mem[1][108] .is_wysiwyg = "true";
defparam \mem[1][108] .power_up = "low";

cyclonev_lcell_comb \mem~11 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][108]~q ),
	.datac(!in_data_reg_108),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~11 .extended_lut = "off";
defparam \mem~11 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~11 .shared_arith = "off";

dffeas \mem[1][109] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][109]~q ),
	.prn(vcc));
defparam \mem[1][109] .is_wysiwyg = "true";
defparam \mem[1][109] .power_up = "low";

cyclonev_lcell_comb \mem~12 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][109]~q ),
	.datac(!in_data_reg_109),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~12 .extended_lut = "off";
defparam \mem~12 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~12 .shared_arith = "off";

dffeas \mem[1][110] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][110]~q ),
	.prn(vcc));
defparam \mem[1][110] .is_wysiwyg = "true";
defparam \mem[1][110] .power_up = "low";

cyclonev_lcell_comb \mem~13 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][110]~q ),
	.datac(!in_data_reg_110),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~13 .extended_lut = "off";
defparam \mem~13 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~13 .shared_arith = "off";

dffeas \mem[1][111] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][111]~q ),
	.prn(vcc));
defparam \mem[1][111] .is_wysiwyg = "true";
defparam \mem[1][111] .power_up = "low";

cyclonev_lcell_comb \mem~14 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][111]~q ),
	.datac(!in_data_reg_111),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~14 .extended_lut = "off";
defparam \mem~14 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~14 .shared_arith = "off";

dffeas \mem[1][112] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][112]~q ),
	.prn(vcc));
defparam \mem[1][112] .is_wysiwyg = "true";
defparam \mem[1][112] .power_up = "low";

cyclonev_lcell_comb \mem~15 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][112]~q ),
	.datac(!in_data_reg_112),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~15 .extended_lut = "off";
defparam \mem~15 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~15 .shared_arith = "off";

dffeas \mem[1][113] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][113]~q ),
	.prn(vcc));
defparam \mem[1][113] .is_wysiwyg = "true";
defparam \mem[1][113] .power_up = "low";

cyclonev_lcell_comb \mem~16 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][113]~q ),
	.datac(!in_data_reg_113),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~16 .extended_lut = "off";
defparam \mem~16 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~16 .shared_arith = "off";

dffeas \mem[1][114] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][114]~q ),
	.prn(vcc));
defparam \mem[1][114] .is_wysiwyg = "true";
defparam \mem[1][114] .power_up = "low";

cyclonev_lcell_comb \mem~17 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][114]~q ),
	.datac(!in_data_reg_114),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~17 .extended_lut = "off";
defparam \mem~17 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~17 .shared_arith = "off";

dffeas \mem[1][115] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][115]~q ),
	.prn(vcc));
defparam \mem[1][115] .is_wysiwyg = "true";
defparam \mem[1][115] .power_up = "low";

cyclonev_lcell_comb \mem~18 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][115]~q ),
	.datac(!in_data_reg_115),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~18 .extended_lut = "off";
defparam \mem~18 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~18 .shared_arith = "off";

dffeas \mem[1][116] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][116]~q ),
	.prn(vcc));
defparam \mem[1][116] .is_wysiwyg = "true";
defparam \mem[1][116] .power_up = "low";

cyclonev_lcell_comb \mem~19 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][116]~q ),
	.datac(!in_data_reg_116),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~19 .extended_lut = "off";
defparam \mem~19 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~19 .shared_arith = "off";

endmodule

module spw_babasu_altera_avalon_sc_fifo_20 (
	read_latency_shift_reg_0,
	mem_used_0,
	mem_129_0,
	mem_used_01,
	av_readdata_pre_0,
	mem_0_0,
	reset,
	WideOr0,
	clk)/* synthesis synthesis_greybox=0 */;
input 	read_latency_shift_reg_0;
output 	mem_used_0;
input 	mem_129_0;
input 	mem_used_01;
input 	av_readdata_pre_0;
output 	mem_0_0;
input 	reset;
input 	WideOr0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~q ;
wire \mem_used[0]~0_combout ;
wire \mem[1][0]~q ;
wire \mem~0_combout ;
wire \mem[0][0]~1_combout ;


dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][0] (
	.clk(clk),
	.d(\mem[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_0_0),
	.prn(vcc));
defparam \mem[0][0] .is_wysiwyg = "true";
defparam \mem[0][0] .power_up = "low";

cyclonev_lcell_comb \read~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_129_0),
	.datad(!mem_used_01),
	.datae(!WideOr0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h0000777000007770;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!\mem_used[1]~q ),
	.datad(!\read~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'h1F001F001F001F00;
defparam \mem_used[1]~1 .shared_arith = "off";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[1]~q ),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!\mem_used[1]~q ),
	.datad(!\read~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~0 .extended_lut = "off";
defparam \mem_used[0]~0 .lut_mask = 64'h731F731F731F731F;
defparam \mem_used[0]~0 .shared_arith = "off";

dffeas \mem[1][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][0]~q ),
	.prn(vcc));
defparam \mem[1][0] .is_wysiwyg = "true";
defparam \mem[1][0] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!av_readdata_pre_0),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h4747474747474747;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \mem[0][0]~1 (
	.dataa(!mem_used_0),
	.datab(!mem_0_0),
	.datac(!\read~0_combout ),
	.datad(!\mem~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem[0][0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem[0][0]~1 .extended_lut = "off";
defparam \mem[0][0]~1 .lut_mask = 64'h10BF10BF10BF10BF;
defparam \mem[0][0]~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_avalon_sc_fifo_21 (
	out_valid_reg,
	mem_used_1,
	WideOr0,
	in_data_reg_68,
	stateST_UNCOMP_WR_SUBBURST,
	mem_129_0,
	mem_used_0,
	mem_68_0,
	mem_66_0,
	comb,
	mem_130_0,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	mem_105_0,
	mem_106_0,
	mem_107_0,
	mem_108_0,
	mem_109_0,
	mem_110_0,
	mem_111_0,
	mem_112_0,
	mem_113_0,
	mem_114_0,
	mem_115_0,
	mem_116_0,
	reset,
	nxt_out_eop,
	last_packet_beat,
	WideOr01,
	read,
	cp_ready,
	in_data_reg_69,
	rf_source_valid,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_6,
	rp_valid,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	clk)/* synthesis synthesis_greybox=0 */;
input 	out_valid_reg;
output 	mem_used_1;
input 	WideOr0;
input 	in_data_reg_68;
input 	stateST_UNCOMP_WR_SUBBURST;
output 	mem_129_0;
output 	mem_used_0;
output 	mem_68_0;
output 	mem_66_0;
input 	comb;
output 	mem_130_0;
output 	mem_78_0;
output 	mem_77_0;
output 	mem_76_0;
output 	mem_75_0;
output 	mem_74_0;
output 	mem_105_0;
output 	mem_106_0;
output 	mem_107_0;
output 	mem_108_0;
output 	mem_109_0;
output 	mem_110_0;
output 	mem_111_0;
output 	mem_112_0;
output 	mem_113_0;
output 	mem_114_0;
output 	mem_115_0;
output 	mem_116_0;
input 	reset;
input 	nxt_out_eop;
input 	last_packet_beat;
input 	WideOr01;
output 	read;
input 	cp_ready;
input 	in_data_reg_69;
input 	rf_source_valid;
input 	out_byte_cnt_reg_2;
input 	out_uncomp_byte_cnt_reg_5;
input 	out_uncomp_byte_cnt_reg_4;
input 	out_uncomp_byte_cnt_reg_3;
input 	out_uncomp_byte_cnt_reg_2;
input 	out_uncomp_byte_cnt_reg_6;
input 	rp_valid;
input 	in_data_reg_105;
input 	in_data_reg_106;
input 	in_data_reg_107;
input 	in_data_reg_108;
input 	in_data_reg_109;
input 	in_data_reg_110;
input 	in_data_reg_111;
input 	in_data_reg_112;
input 	in_data_reg_113;
input 	in_data_reg_114;
input 	in_data_reg_115;
input 	in_data_reg_116;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \write~0_combout ;
wire \mem_used[1]~0_combout ;
wire \mem[1][129]~q ;
wire \mem~20_combout ;
wire \always0~0_combout ;
wire \mem_used[0]~1_combout ;
wire \mem[1][68]~q ;
wire \mem~0_combout ;
wire \mem[1][69]~q ;
wire \mem~1_combout ;
wire \mem[1][130]~q ;
wire \mem~2_combout ;
wire \mem[1][78]~q ;
wire \mem~3_combout ;
wire \mem[1][77]~q ;
wire \mem~4_combout ;
wire \mem[1][76]~q ;
wire \mem~5_combout ;
wire \mem[1][75]~q ;
wire \mem~6_combout ;
wire \mem[1][74]~q ;
wire \mem~7_combout ;
wire \mem[1][105]~q ;
wire \mem~8_combout ;
wire \mem[1][106]~q ;
wire \mem~9_combout ;
wire \mem[1][107]~q ;
wire \mem~10_combout ;
wire \mem[1][108]~q ;
wire \mem~11_combout ;
wire \mem[1][109]~q ;
wire \mem~12_combout ;
wire \mem[1][110]~q ;
wire \mem~13_combout ;
wire \mem[1][111]~q ;
wire \mem~14_combout ;
wire \mem[1][112]~q ;
wire \mem~15_combout ;
wire \mem[1][113]~q ;
wire \mem~16_combout ;
wire \mem[1][114]~q ;
wire \mem~17_combout ;
wire \mem[1][115]~q ;
wire \mem~18_combout ;
wire \mem[1][116]~q ;
wire \mem~19_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][129] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_129_0),
	.prn(vcc));
defparam \mem[0][129] .is_wysiwyg = "true";
defparam \mem[0][129] .power_up = "low";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][68] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_68_0),
	.prn(vcc));
defparam \mem[0][68] .is_wysiwyg = "true";
defparam \mem[0][68] .power_up = "low";

dffeas \mem[0][66] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_66_0),
	.prn(vcc));
defparam \mem[0][66] .is_wysiwyg = "true";
defparam \mem[0][66] .power_up = "low";

dffeas \mem[0][130] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_130_0),
	.prn(vcc));
defparam \mem[0][130] .is_wysiwyg = "true";
defparam \mem[0][130] .power_up = "low";

dffeas \mem[0][78] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_78_0),
	.prn(vcc));
defparam \mem[0][78] .is_wysiwyg = "true";
defparam \mem[0][78] .power_up = "low";

dffeas \mem[0][77] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_77_0),
	.prn(vcc));
defparam \mem[0][77] .is_wysiwyg = "true";
defparam \mem[0][77] .power_up = "low";

dffeas \mem[0][76] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_76_0),
	.prn(vcc));
defparam \mem[0][76] .is_wysiwyg = "true";
defparam \mem[0][76] .power_up = "low";

dffeas \mem[0][75] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_75_0),
	.prn(vcc));
defparam \mem[0][75] .is_wysiwyg = "true";
defparam \mem[0][75] .power_up = "low";

dffeas \mem[0][74] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_74_0),
	.prn(vcc));
defparam \mem[0][74] .is_wysiwyg = "true";
defparam \mem[0][74] .power_up = "low";

dffeas \mem[0][105] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_105_0),
	.prn(vcc));
defparam \mem[0][105] .is_wysiwyg = "true";
defparam \mem[0][105] .power_up = "low";

dffeas \mem[0][106] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_106_0),
	.prn(vcc));
defparam \mem[0][106] .is_wysiwyg = "true";
defparam \mem[0][106] .power_up = "low";

dffeas \mem[0][107] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_107_0),
	.prn(vcc));
defparam \mem[0][107] .is_wysiwyg = "true";
defparam \mem[0][107] .power_up = "low";

dffeas \mem[0][108] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_108_0),
	.prn(vcc));
defparam \mem[0][108] .is_wysiwyg = "true";
defparam \mem[0][108] .power_up = "low";

dffeas \mem[0][109] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_109_0),
	.prn(vcc));
defparam \mem[0][109] .is_wysiwyg = "true";
defparam \mem[0][109] .power_up = "low";

dffeas \mem[0][110] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_110_0),
	.prn(vcc));
defparam \mem[0][110] .is_wysiwyg = "true";
defparam \mem[0][110] .power_up = "low";

dffeas \mem[0][111] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_111_0),
	.prn(vcc));
defparam \mem[0][111] .is_wysiwyg = "true";
defparam \mem[0][111] .power_up = "low";

dffeas \mem[0][112] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_112_0),
	.prn(vcc));
defparam \mem[0][112] .is_wysiwyg = "true";
defparam \mem[0][112] .power_up = "low";

dffeas \mem[0][113] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_113_0),
	.prn(vcc));
defparam \mem[0][113] .is_wysiwyg = "true";
defparam \mem[0][113] .power_up = "low";

dffeas \mem[0][114] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_114_0),
	.prn(vcc));
defparam \mem[0][114] .is_wysiwyg = "true";
defparam \mem[0][114] .power_up = "low";

dffeas \mem[0][115] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_115_0),
	.prn(vcc));
defparam \mem[0][115] .is_wysiwyg = "true";
defparam \mem[0][115] .power_up = "low";

dffeas \mem[0][116] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_116_0),
	.prn(vcc));
defparam \mem[0][116] .is_wysiwyg = "true";
defparam \mem[0][116] .power_up = "low";

cyclonev_lcell_comb \read~0 (
	.dataa(!comb),
	.datab(!WideOr01),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h1111111111111111;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \write~0 (
	.dataa(!mem_used_1),
	.datab(!WideOr0),
	.datac(!cp_ready),
	.datad(!rf_source_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'h008A008A008A008A;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!last_packet_beat),
	.datad(!read),
	.datae(!\write~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'h5505335355053353;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][129] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][129]~q ),
	.prn(vcc));
defparam \mem[1][129] .is_wysiwyg = "true";
defparam \mem[1][129] .power_up = "low";

cyclonev_lcell_comb \mem~20 (
	.dataa(!WideOr0),
	.datab(!out_valid_reg),
	.datac(!\mem[1][129]~q ),
	.datad(!in_data_reg_68),
	.datae(!mem_used_1),
	.dataf(!nxt_out_eop),
	.datag(!in_data_reg_69),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~20 .extended_lut = "on";
defparam \mem~20 .lut_mask = 64'h02020F0F02330F0F;
defparam \mem~20 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!mem_used_0),
	.datab(!rp_valid),
	.datac(!last_packet_beat),
	.datad(!read),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hAAEAAAEAAAEAAAEA;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!rp_valid),
	.datad(!last_packet_beat),
	.datae(!read),
	.dataf(!\write~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'h33331333FFFFFFFF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem[1][68] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][68]~q ),
	.prn(vcc));
defparam \mem[1][68] .is_wysiwyg = "true";
defparam \mem[1][68] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!mem_used_1),
	.datab(!in_data_reg_68),
	.datac(!\mem[1][68]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h2727272727272727;
defparam \mem~0 .shared_arith = "off";

dffeas \mem[1][69] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][69]~q ),
	.prn(vcc));
defparam \mem[1][69] .is_wysiwyg = "true";
defparam \mem[1][69] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!mem_used_1),
	.datab(!in_data_reg_69),
	.datac(!\mem[1][69]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h2727272727272727;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[1][130] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][130]~q ),
	.prn(vcc));
defparam \mem[1][130] .is_wysiwyg = "true";
defparam \mem[1][130] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!mem_used_1),
	.datab(!nxt_out_eop),
	.datac(!\mem[1][130]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h2727272727272727;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[1][78] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][78]~q ),
	.prn(vcc));
defparam \mem[1][78] .is_wysiwyg = "true";
defparam \mem[1][78] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_6),
	.datad(!\mem[1][78]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h0257025702570257;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][77] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][77]~q ),
	.prn(vcc));
defparam \mem[1][77] .is_wysiwyg = "true";
defparam \mem[1][77] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\mem[1][77]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h0257025702570257;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][76] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][76]~q ),
	.prn(vcc));
defparam \mem[1][76] .is_wysiwyg = "true";
defparam \mem[1][76] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!\mem[1][76]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h0257025702570257;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][75] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][75]~q ),
	.prn(vcc));
defparam \mem[1][75] .is_wysiwyg = "true";
defparam \mem[1][75] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\mem[1][75]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h0257025702570257;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[1][74] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][74]~q ),
	.prn(vcc));
defparam \mem[1][74] .is_wysiwyg = "true";
defparam \mem[1][74] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_byte_cnt_reg_2),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(!\mem[1][74]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h082A5D7F082A5D7F;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[1][105] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][105]~q ),
	.prn(vcc));
defparam \mem[1][105] .is_wysiwyg = "true";
defparam \mem[1][105] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][105]~q ),
	.datac(!in_data_reg_105),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~8 .shared_arith = "off";

dffeas \mem[1][106] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][106]~q ),
	.prn(vcc));
defparam \mem[1][106] .is_wysiwyg = "true";
defparam \mem[1][106] .power_up = "low";

cyclonev_lcell_comb \mem~9 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][106]~q ),
	.datac(!in_data_reg_106),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~9 .extended_lut = "off";
defparam \mem~9 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~9 .shared_arith = "off";

dffeas \mem[1][107] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][107]~q ),
	.prn(vcc));
defparam \mem[1][107] .is_wysiwyg = "true";
defparam \mem[1][107] .power_up = "low";

cyclonev_lcell_comb \mem~10 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][107]~q ),
	.datac(!in_data_reg_107),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~10 .extended_lut = "off";
defparam \mem~10 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~10 .shared_arith = "off";

dffeas \mem[1][108] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][108]~q ),
	.prn(vcc));
defparam \mem[1][108] .is_wysiwyg = "true";
defparam \mem[1][108] .power_up = "low";

cyclonev_lcell_comb \mem~11 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][108]~q ),
	.datac(!in_data_reg_108),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~11 .extended_lut = "off";
defparam \mem~11 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~11 .shared_arith = "off";

dffeas \mem[1][109] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][109]~q ),
	.prn(vcc));
defparam \mem[1][109] .is_wysiwyg = "true";
defparam \mem[1][109] .power_up = "low";

cyclonev_lcell_comb \mem~12 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][109]~q ),
	.datac(!in_data_reg_109),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~12 .extended_lut = "off";
defparam \mem~12 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~12 .shared_arith = "off";

dffeas \mem[1][110] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][110]~q ),
	.prn(vcc));
defparam \mem[1][110] .is_wysiwyg = "true";
defparam \mem[1][110] .power_up = "low";

cyclonev_lcell_comb \mem~13 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][110]~q ),
	.datac(!in_data_reg_110),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~13 .extended_lut = "off";
defparam \mem~13 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~13 .shared_arith = "off";

dffeas \mem[1][111] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][111]~q ),
	.prn(vcc));
defparam \mem[1][111] .is_wysiwyg = "true";
defparam \mem[1][111] .power_up = "low";

cyclonev_lcell_comb \mem~14 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][111]~q ),
	.datac(!in_data_reg_111),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~14 .extended_lut = "off";
defparam \mem~14 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~14 .shared_arith = "off";

dffeas \mem[1][112] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][112]~q ),
	.prn(vcc));
defparam \mem[1][112] .is_wysiwyg = "true";
defparam \mem[1][112] .power_up = "low";

cyclonev_lcell_comb \mem~15 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][112]~q ),
	.datac(!in_data_reg_112),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~15 .extended_lut = "off";
defparam \mem~15 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~15 .shared_arith = "off";

dffeas \mem[1][113] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][113]~q ),
	.prn(vcc));
defparam \mem[1][113] .is_wysiwyg = "true";
defparam \mem[1][113] .power_up = "low";

cyclonev_lcell_comb \mem~16 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][113]~q ),
	.datac(!in_data_reg_113),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~16 .extended_lut = "off";
defparam \mem~16 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~16 .shared_arith = "off";

dffeas \mem[1][114] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][114]~q ),
	.prn(vcc));
defparam \mem[1][114] .is_wysiwyg = "true";
defparam \mem[1][114] .power_up = "low";

cyclonev_lcell_comb \mem~17 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][114]~q ),
	.datac(!in_data_reg_114),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~17 .extended_lut = "off";
defparam \mem~17 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~17 .shared_arith = "off";

dffeas \mem[1][115] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][115]~q ),
	.prn(vcc));
defparam \mem[1][115] .is_wysiwyg = "true";
defparam \mem[1][115] .power_up = "low";

cyclonev_lcell_comb \mem~18 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][115]~q ),
	.datac(!in_data_reg_115),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~18 .extended_lut = "off";
defparam \mem~18 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~18 .shared_arith = "off";

dffeas \mem[1][116] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][116]~q ),
	.prn(vcc));
defparam \mem[1][116] .is_wysiwyg = "true";
defparam \mem[1][116] .power_up = "low";

cyclonev_lcell_comb \mem~19 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][116]~q ),
	.datac(!in_data_reg_116),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~19 .extended_lut = "off";
defparam \mem~19 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~19 .shared_arith = "off";

endmodule

module spw_babasu_altera_avalon_sc_fifo_22 (
	h2f_RREADY_0,
	read_latency_shift_reg_0,
	mem_used_0,
	empty1,
	av_readdata_pre_0,
	mem_0_0,
	reset,
	clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_RREADY_0;
input 	read_latency_shift_reg_0;
output 	mem_used_0;
output 	empty1;
input 	av_readdata_pre_0;
output 	mem_0_0;
input 	reset;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[1]~1_combout ;
wire \mem_used[1]~q ;
wire \mem_used[0]~0_combout ;
wire \mem[1][0]~q ;
wire \mem~0_combout ;
wire \mem[0][0]~1_combout ;


dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb empty(
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(empty1),
	.sumout(),
	.cout(),
	.shareout());
defparam empty.extended_lut = "off";
defparam empty.lut_mask = 64'h8888888888888888;
defparam empty.shared_arith = "off";

dffeas \mem[0][0] (
	.clk(clk),
	.d(\mem[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_0_0),
	.prn(vcc));
defparam \mem[0][0] .is_wysiwyg = "true";
defparam \mem[0][0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!h2f_RREADY_0),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem_used[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'h02EA02EA02EA02EA;
defparam \mem_used[1]~1 .shared_arith = "off";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[1]~q ),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~0 (
	.dataa(!h2f_RREADY_0),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem_used[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~0 .extended_lut = "off";
defparam \mem_used[0]~0 .lut_mask = 64'h2B1F2B1F2B1F2B1F;
defparam \mem_used[0]~0 .shared_arith = "off";

dffeas \mem[1][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][0]~q ),
	.prn(vcc));
defparam \mem[1][0] .is_wysiwyg = "true";
defparam \mem[1][0] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!av_readdata_pre_0),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h4747474747474747;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \mem[0][0]~1 (
	.dataa(!h2f_RREADY_0),
	.datab(!mem_used_0),
	.datac(!mem_0_0),
	.datad(!\mem~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem[0][0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem[0][0]~1 .extended_lut = "off";
defparam \mem[0][0]~1 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \mem[0][0]~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_avalon_sc_fifo_23 (
	h2f_RREADY_0,
	waitrequest_reset_override,
	mem_used_1,
	in_data_reg_69,
	wait_latency_counter_1,
	wait_latency_counter_0,
	nxt_out_eop,
	out_valid_reg,
	stateST_UNCOMP_WR_SUBBURST,
	mem_130_0,
	empty,
	mem_66_0,
	mem_used_0,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	mem_105_0,
	mem_106_0,
	mem_107_0,
	mem_108_0,
	mem_109_0,
	mem_110_0,
	mem_111_0,
	mem_112_0,
	mem_113_0,
	mem_114_0,
	mem_115_0,
	mem_116_0,
	reset,
	last_packet_beat,
	write,
	write1,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_6,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_RREADY_0;
input 	waitrequest_reset_override;
output 	mem_used_1;
input 	in_data_reg_69;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	nxt_out_eop;
input 	out_valid_reg;
input 	stateST_UNCOMP_WR_SUBBURST;
output 	mem_130_0;
input 	empty;
output 	mem_66_0;
output 	mem_used_0;
output 	mem_78_0;
output 	mem_77_0;
output 	mem_76_0;
output 	mem_75_0;
output 	mem_74_0;
output 	mem_105_0;
output 	mem_106_0;
output 	mem_107_0;
output 	mem_108_0;
output 	mem_109_0;
output 	mem_110_0;
output 	mem_111_0;
output 	mem_112_0;
output 	mem_113_0;
output 	mem_114_0;
output 	mem_115_0;
output 	mem_116_0;
input 	reset;
input 	last_packet_beat;
output 	write;
output 	write1;
input 	out_byte_cnt_reg_2;
input 	out_uncomp_byte_cnt_reg_3;
input 	out_uncomp_byte_cnt_reg_2;
input 	out_uncomp_byte_cnt_reg_4;
input 	out_uncomp_byte_cnt_reg_5;
input 	out_uncomp_byte_cnt_reg_6;
input 	in_data_reg_105;
input 	in_data_reg_106;
input 	in_data_reg_107;
input 	in_data_reg_108;
input 	in_data_reg_109;
input 	in_data_reg_110;
input 	in_data_reg_111;
input 	in_data_reg_112;
input 	in_data_reg_113;
input 	in_data_reg_114;
input 	in_data_reg_115;
input 	in_data_reg_116;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read~0_combout ;
wire \mem_used[1]~0_combout ;
wire \mem[1][130]~q ;
wire \mem~0_combout ;
wire \always0~0_combout ;
wire \mem[1][69]~q ;
wire \mem~1_combout ;
wire \mem_used[0]~1_combout ;
wire \mem[1][78]~q ;
wire \mem~2_combout ;
wire \mem[1][77]~q ;
wire \mem~3_combout ;
wire \mem[1][76]~q ;
wire \mem~4_combout ;
wire \mem[1][75]~q ;
wire \mem~5_combout ;
wire \mem[1][74]~q ;
wire \mem~6_combout ;
wire \mem[1][105]~q ;
wire \mem~7_combout ;
wire \mem[1][106]~q ;
wire \mem~8_combout ;
wire \mem[1][107]~q ;
wire \mem~9_combout ;
wire \mem[1][108]~q ;
wire \mem~10_combout ;
wire \mem[1][109]~q ;
wire \mem~11_combout ;
wire \mem[1][110]~q ;
wire \mem~12_combout ;
wire \mem[1][111]~q ;
wire \mem~13_combout ;
wire \mem[1][112]~q ;
wire \mem~14_combout ;
wire \mem[1][113]~q ;
wire \mem~15_combout ;
wire \mem[1][114]~q ;
wire \mem~16_combout ;
wire \mem[1][115]~q ;
wire \mem~17_combout ;
wire \mem[1][116]~q ;
wire \mem~18_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][130] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_130_0),
	.prn(vcc));
defparam \mem[0][130] .is_wysiwyg = "true";
defparam \mem[0][130] .power_up = "low";

dffeas \mem[0][66] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_66_0),
	.prn(vcc));
defparam \mem[0][66] .is_wysiwyg = "true";
defparam \mem[0][66] .power_up = "low";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][78] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_78_0),
	.prn(vcc));
defparam \mem[0][78] .is_wysiwyg = "true";
defparam \mem[0][78] .power_up = "low";

dffeas \mem[0][77] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_77_0),
	.prn(vcc));
defparam \mem[0][77] .is_wysiwyg = "true";
defparam \mem[0][77] .power_up = "low";

dffeas \mem[0][76] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_76_0),
	.prn(vcc));
defparam \mem[0][76] .is_wysiwyg = "true";
defparam \mem[0][76] .power_up = "low";

dffeas \mem[0][75] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_75_0),
	.prn(vcc));
defparam \mem[0][75] .is_wysiwyg = "true";
defparam \mem[0][75] .power_up = "low";

dffeas \mem[0][74] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_74_0),
	.prn(vcc));
defparam \mem[0][74] .is_wysiwyg = "true";
defparam \mem[0][74] .power_up = "low";

dffeas \mem[0][105] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_105_0),
	.prn(vcc));
defparam \mem[0][105] .is_wysiwyg = "true";
defparam \mem[0][105] .power_up = "low";

dffeas \mem[0][106] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_106_0),
	.prn(vcc));
defparam \mem[0][106] .is_wysiwyg = "true";
defparam \mem[0][106] .power_up = "low";

dffeas \mem[0][107] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_107_0),
	.prn(vcc));
defparam \mem[0][107] .is_wysiwyg = "true";
defparam \mem[0][107] .power_up = "low";

dffeas \mem[0][108] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_108_0),
	.prn(vcc));
defparam \mem[0][108] .is_wysiwyg = "true";
defparam \mem[0][108] .power_up = "low";

dffeas \mem[0][109] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_109_0),
	.prn(vcc));
defparam \mem[0][109] .is_wysiwyg = "true";
defparam \mem[0][109] .power_up = "low";

dffeas \mem[0][110] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_110_0),
	.prn(vcc));
defparam \mem[0][110] .is_wysiwyg = "true";
defparam \mem[0][110] .power_up = "low";

dffeas \mem[0][111] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_111_0),
	.prn(vcc));
defparam \mem[0][111] .is_wysiwyg = "true";
defparam \mem[0][111] .power_up = "low";

dffeas \mem[0][112] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_112_0),
	.prn(vcc));
defparam \mem[0][112] .is_wysiwyg = "true";
defparam \mem[0][112] .power_up = "low";

dffeas \mem[0][113] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_113_0),
	.prn(vcc));
defparam \mem[0][113] .is_wysiwyg = "true";
defparam \mem[0][113] .power_up = "low";

dffeas \mem[0][114] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_114_0),
	.prn(vcc));
defparam \mem[0][114] .is_wysiwyg = "true";
defparam \mem[0][114] .power_up = "low";

dffeas \mem[0][115] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_115_0),
	.prn(vcc));
defparam \mem[0][115] .is_wysiwyg = "true";
defparam \mem[0][115] .power_up = "low";

dffeas \mem[0][116] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_116_0),
	.prn(vcc));
defparam \mem[0][116] .is_wysiwyg = "true";
defparam \mem[0][116] .power_up = "low";

cyclonev_lcell_comb \write~0 (
	.dataa(!waitrequest_reset_override),
	.datab(!in_data_reg_69),
	.datac(!mem_used_1),
	.datad(!out_valid_reg),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'h0010001000100010;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \write~1 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!write),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write1),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~1 .extended_lut = "off";
defparam \write~1 .lut_mask = 64'h0202020202020202;
defparam \write~1 .shared_arith = "off";

cyclonev_lcell_comb \read~0 (
	.dataa(!h2f_RREADY_0),
	.datab(!empty),
	.datac(!last_packet_beat),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h4040404040404040;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!\read~0_combout ),
	.datad(!write1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'h5431543154315431;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][130] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][130]~q ),
	.prn(vcc));
defparam \mem[1][130] .is_wysiwyg = "true";
defparam \mem[1][130] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!mem_used_1),
	.datab(!nxt_out_eop),
	.datac(!\mem[1][130]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h2727272727272727;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!mem_used_0),
	.datab(!\read~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \always0~0 .shared_arith = "off";

dffeas \mem[1][69] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][69]~q ),
	.prn(vcc));
defparam \mem[1][69] .is_wysiwyg = "true";
defparam \mem[1][69] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!in_data_reg_69),
	.datab(!mem_used_1),
	.datac(!\mem[1][69]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h4747474747474747;
defparam \mem~1 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!\read~0_combout ),
	.datad(!write1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'h31FF31FF31FF31FF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem[1][78] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][78]~q ),
	.prn(vcc));
defparam \mem[1][78] .is_wysiwyg = "true";
defparam \mem[1][78] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_6),
	.datad(!\mem[1][78]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h0257025702570257;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[1][77] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][77]~q ),
	.prn(vcc));
defparam \mem[1][77] .is_wysiwyg = "true";
defparam \mem[1][77] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\mem[1][77]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h0257025702570257;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][76] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][76]~q ),
	.prn(vcc));
defparam \mem[1][76] .is_wysiwyg = "true";
defparam \mem[1][76] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!\mem[1][76]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h0257025702570257;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][75] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][75]~q ),
	.prn(vcc));
defparam \mem[1][75] .is_wysiwyg = "true";
defparam \mem[1][75] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\mem[1][75]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h0257025702570257;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][74] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][74]~q ),
	.prn(vcc));
defparam \mem[1][74] .is_wysiwyg = "true";
defparam \mem[1][74] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_byte_cnt_reg_2),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(!\mem[1][74]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h082A5D7F082A5D7F;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[1][105] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][105]~q ),
	.prn(vcc));
defparam \mem[1][105] .is_wysiwyg = "true";
defparam \mem[1][105] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][105]~q ),
	.datac(!in_data_reg_105),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[1][106] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][106]~q ),
	.prn(vcc));
defparam \mem[1][106] .is_wysiwyg = "true";
defparam \mem[1][106] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][106]~q ),
	.datac(!in_data_reg_106),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~8 .shared_arith = "off";

dffeas \mem[1][107] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][107]~q ),
	.prn(vcc));
defparam \mem[1][107] .is_wysiwyg = "true";
defparam \mem[1][107] .power_up = "low";

cyclonev_lcell_comb \mem~9 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][107]~q ),
	.datac(!in_data_reg_107),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~9 .extended_lut = "off";
defparam \mem~9 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~9 .shared_arith = "off";

dffeas \mem[1][108] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][108]~q ),
	.prn(vcc));
defparam \mem[1][108] .is_wysiwyg = "true";
defparam \mem[1][108] .power_up = "low";

cyclonev_lcell_comb \mem~10 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][108]~q ),
	.datac(!in_data_reg_108),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~10 .extended_lut = "off";
defparam \mem~10 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~10 .shared_arith = "off";

dffeas \mem[1][109] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][109]~q ),
	.prn(vcc));
defparam \mem[1][109] .is_wysiwyg = "true";
defparam \mem[1][109] .power_up = "low";

cyclonev_lcell_comb \mem~11 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][109]~q ),
	.datac(!in_data_reg_109),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~11 .extended_lut = "off";
defparam \mem~11 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~11 .shared_arith = "off";

dffeas \mem[1][110] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][110]~q ),
	.prn(vcc));
defparam \mem[1][110] .is_wysiwyg = "true";
defparam \mem[1][110] .power_up = "low";

cyclonev_lcell_comb \mem~12 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][110]~q ),
	.datac(!in_data_reg_110),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~12 .extended_lut = "off";
defparam \mem~12 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~12 .shared_arith = "off";

dffeas \mem[1][111] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][111]~q ),
	.prn(vcc));
defparam \mem[1][111] .is_wysiwyg = "true";
defparam \mem[1][111] .power_up = "low";

cyclonev_lcell_comb \mem~13 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][111]~q ),
	.datac(!in_data_reg_111),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~13 .extended_lut = "off";
defparam \mem~13 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~13 .shared_arith = "off";

dffeas \mem[1][112] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][112]~q ),
	.prn(vcc));
defparam \mem[1][112] .is_wysiwyg = "true";
defparam \mem[1][112] .power_up = "low";

cyclonev_lcell_comb \mem~14 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][112]~q ),
	.datac(!in_data_reg_112),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~14 .extended_lut = "off";
defparam \mem~14 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~14 .shared_arith = "off";

dffeas \mem[1][113] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][113]~q ),
	.prn(vcc));
defparam \mem[1][113] .is_wysiwyg = "true";
defparam \mem[1][113] .power_up = "low";

cyclonev_lcell_comb \mem~15 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][113]~q ),
	.datac(!in_data_reg_113),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~15 .extended_lut = "off";
defparam \mem~15 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~15 .shared_arith = "off";

dffeas \mem[1][114] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][114]~q ),
	.prn(vcc));
defparam \mem[1][114] .is_wysiwyg = "true";
defparam \mem[1][114] .power_up = "low";

cyclonev_lcell_comb \mem~16 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][114]~q ),
	.datac(!in_data_reg_114),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~16 .extended_lut = "off";
defparam \mem~16 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~16 .shared_arith = "off";

dffeas \mem[1][115] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][115]~q ),
	.prn(vcc));
defparam \mem[1][115] .is_wysiwyg = "true";
defparam \mem[1][115] .power_up = "low";

cyclonev_lcell_comb \mem~17 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][115]~q ),
	.datac(!in_data_reg_115),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~17 .extended_lut = "off";
defparam \mem~17 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~17 .shared_arith = "off";

dffeas \mem[1][116] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][116]~q ),
	.prn(vcc));
defparam \mem[1][116] .is_wysiwyg = "true";
defparam \mem[1][116] .power_up = "low";

cyclonev_lcell_comb \mem~18 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][116]~q ),
	.datac(!in_data_reg_116),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~18 .extended_lut = "off";
defparam \mem~18 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~18 .shared_arith = "off";

endmodule

module spw_babasu_altera_avalon_sc_fifo_24 (
	read_latency_shift_reg_0,
	mem_used_0,
	mem_129_0,
	mem_used_01,
	av_readdata_pre_0,
	always4,
	mem_0_0,
	av_readdata_pre_1,
	mem_1_0,
	av_readdata_pre_2,
	mem_2_0,
	av_readdata_pre_3,
	mem_3_0,
	av_readdata_pre_4,
	mem_4_0,
	av_readdata_pre_5,
	mem_5_0,
	av_readdata_pre_6,
	mem_6_0,
	av_readdata_pre_7,
	mem_7_0,
	reset,
	WideOr0,
	clk)/* synthesis synthesis_greybox=0 */;
input 	read_latency_shift_reg_0;
output 	mem_used_0;
input 	mem_129_0;
input 	mem_used_01;
input 	av_readdata_pre_0;
output 	always4;
output 	mem_0_0;
input 	av_readdata_pre_1;
output 	mem_1_0;
input 	av_readdata_pre_2;
output 	mem_2_0;
input 	av_readdata_pre_3;
output 	mem_3_0;
input 	av_readdata_pre_4;
output 	mem_4_0;
input 	av_readdata_pre_5;
output 	mem_5_0;
input 	av_readdata_pre_6;
output 	mem_6_0;
input 	av_readdata_pre_7;
output 	mem_7_0;
input 	reset;
input 	WideOr0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~q ;
wire \mem_used[0]~0_combout ;
wire \mem[1][0]~q ;
wire \mem~0_combout ;
wire \always0~0_combout ;
wire \mem[1][1]~q ;
wire \mem~1_combout ;
wire \mem[1][2]~q ;
wire \mem~2_combout ;
wire \mem[1][3]~q ;
wire \mem~3_combout ;
wire \mem[1][4]~q ;
wire \mem~4_combout ;
wire \mem[1][5]~q ;
wire \mem~5_combout ;
wire \mem[1][6]~q ;
wire \mem~6_combout ;
wire \mem[1][7]~q ;
wire \mem~7_combout ;


dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \always4~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always4),
	.sumout(),
	.cout(),
	.shareout());
defparam \always4~0 .extended_lut = "off";
defparam \always4~0 .lut_mask = 64'h4444444444444444;
defparam \always4~0 .shared_arith = "off";

dffeas \mem[0][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_0_0),
	.prn(vcc));
defparam \mem[0][0] .is_wysiwyg = "true";
defparam \mem[0][0] .power_up = "low";

dffeas \mem[0][1] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_1_0),
	.prn(vcc));
defparam \mem[0][1] .is_wysiwyg = "true";
defparam \mem[0][1] .power_up = "low";

dffeas \mem[0][2] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_2_0),
	.prn(vcc));
defparam \mem[0][2] .is_wysiwyg = "true";
defparam \mem[0][2] .power_up = "low";

dffeas \mem[0][3] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_3_0),
	.prn(vcc));
defparam \mem[0][3] .is_wysiwyg = "true";
defparam \mem[0][3] .power_up = "low";

dffeas \mem[0][4] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_4_0),
	.prn(vcc));
defparam \mem[0][4] .is_wysiwyg = "true";
defparam \mem[0][4] .power_up = "low";

dffeas \mem[0][5] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_5_0),
	.prn(vcc));
defparam \mem[0][5] .is_wysiwyg = "true";
defparam \mem[0][5] .power_up = "low";

dffeas \mem[0][6] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_6_0),
	.prn(vcc));
defparam \mem[0][6] .is_wysiwyg = "true";
defparam \mem[0][6] .power_up = "low";

dffeas \mem[0][7] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_7_0),
	.prn(vcc));
defparam \mem[0][7] .is_wysiwyg = "true";
defparam \mem[0][7] .power_up = "low";

cyclonev_lcell_comb \read~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_129_0),
	.datad(!mem_used_01),
	.datae(!WideOr0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h0000777000007770;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!\mem_used[1]~q ),
	.datad(!\read~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'h1F001F001F001F00;
defparam \mem_used[1]~1 .shared_arith = "off";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[1]~q ),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!\mem_used[1]~q ),
	.datad(!\read~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~0 .extended_lut = "off";
defparam \mem_used[0]~0 .lut_mask = 64'h731F731F731F731F;
defparam \mem_used[0]~0 .shared_arith = "off";

dffeas \mem[1][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][0]~q ),
	.prn(vcc));
defparam \mem[1][0] .is_wysiwyg = "true";
defparam \mem[1][0] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!av_readdata_pre_0),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h4747474747474747;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!mem_used_0),
	.datab(!\read~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \always0~0 .shared_arith = "off";

dffeas \mem[1][1] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][1]~q ),
	.prn(vcc));
defparam \mem[1][1] .is_wysiwyg = "true";
defparam \mem[1][1] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!av_readdata_pre_1),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h4747474747474747;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[1][2] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][2]~q ),
	.prn(vcc));
defparam \mem[1][2] .is_wysiwyg = "true";
defparam \mem[1][2] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!av_readdata_pre_2),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h4747474747474747;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[1][3] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][3]~q ),
	.prn(vcc));
defparam \mem[1][3] .is_wysiwyg = "true";
defparam \mem[1][3] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!av_readdata_pre_3),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h4747474747474747;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][4] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][4]~q ),
	.prn(vcc));
defparam \mem[1][4] .is_wysiwyg = "true";
defparam \mem[1][4] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!av_readdata_pre_4),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h4747474747474747;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][5] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][5]~q ),
	.prn(vcc));
defparam \mem[1][5] .is_wysiwyg = "true";
defparam \mem[1][5] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!av_readdata_pre_5),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][5]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h4747474747474747;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][6] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][6]~q ),
	.prn(vcc));
defparam \mem[1][6] .is_wysiwyg = "true";
defparam \mem[1][6] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!av_readdata_pre_6),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][6]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h4747474747474747;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[1][7] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][7]~q ),
	.prn(vcc));
defparam \mem[1][7] .is_wysiwyg = "true";
defparam \mem[1][7] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!av_readdata_pre_7),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h4747474747474747;
defparam \mem~7 .shared_arith = "off";

endmodule

module spw_babasu_altera_avalon_sc_fifo_25 (
	out_valid_reg,
	mem_used_1,
	WideOr0,
	in_data_reg_68,
	stateST_UNCOMP_WR_SUBBURST,
	mem_129_0,
	mem_used_0,
	mem_68_0,
	mem_66_0,
	comb,
	mem_130_0,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	mem_105_0,
	mem_106_0,
	mem_107_0,
	mem_108_0,
	mem_109_0,
	mem_110_0,
	mem_111_0,
	mem_112_0,
	mem_113_0,
	mem_114_0,
	mem_115_0,
	mem_116_0,
	reset,
	nxt_out_eop,
	last_packet_beat,
	WideOr01,
	read,
	cp_ready,
	in_data_reg_69,
	rf_source_valid,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_6,
	rp_valid,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	clk)/* synthesis synthesis_greybox=0 */;
input 	out_valid_reg;
output 	mem_used_1;
input 	WideOr0;
input 	in_data_reg_68;
input 	stateST_UNCOMP_WR_SUBBURST;
output 	mem_129_0;
output 	mem_used_0;
output 	mem_68_0;
output 	mem_66_0;
input 	comb;
output 	mem_130_0;
output 	mem_78_0;
output 	mem_77_0;
output 	mem_76_0;
output 	mem_75_0;
output 	mem_74_0;
output 	mem_105_0;
output 	mem_106_0;
output 	mem_107_0;
output 	mem_108_0;
output 	mem_109_0;
output 	mem_110_0;
output 	mem_111_0;
output 	mem_112_0;
output 	mem_113_0;
output 	mem_114_0;
output 	mem_115_0;
output 	mem_116_0;
input 	reset;
input 	nxt_out_eop;
input 	last_packet_beat;
input 	WideOr01;
output 	read;
input 	cp_ready;
input 	in_data_reg_69;
input 	rf_source_valid;
input 	out_byte_cnt_reg_2;
input 	out_uncomp_byte_cnt_reg_5;
input 	out_uncomp_byte_cnt_reg_4;
input 	out_uncomp_byte_cnt_reg_3;
input 	out_uncomp_byte_cnt_reg_2;
input 	out_uncomp_byte_cnt_reg_6;
input 	rp_valid;
input 	in_data_reg_105;
input 	in_data_reg_106;
input 	in_data_reg_107;
input 	in_data_reg_108;
input 	in_data_reg_109;
input 	in_data_reg_110;
input 	in_data_reg_111;
input 	in_data_reg_112;
input 	in_data_reg_113;
input 	in_data_reg_114;
input 	in_data_reg_115;
input 	in_data_reg_116;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \write~0_combout ;
wire \mem_used[1]~0_combout ;
wire \mem[1][129]~q ;
wire \mem~20_combout ;
wire \always0~0_combout ;
wire \mem_used[0]~1_combout ;
wire \mem[1][68]~q ;
wire \mem~0_combout ;
wire \mem[1][69]~q ;
wire \mem~1_combout ;
wire \mem[1][130]~q ;
wire \mem~2_combout ;
wire \mem[1][78]~q ;
wire \mem~3_combout ;
wire \mem[1][77]~q ;
wire \mem~4_combout ;
wire \mem[1][76]~q ;
wire \mem~5_combout ;
wire \mem[1][75]~q ;
wire \mem~6_combout ;
wire \mem[1][74]~q ;
wire \mem~7_combout ;
wire \mem[1][105]~q ;
wire \mem~8_combout ;
wire \mem[1][106]~q ;
wire \mem~9_combout ;
wire \mem[1][107]~q ;
wire \mem~10_combout ;
wire \mem[1][108]~q ;
wire \mem~11_combout ;
wire \mem[1][109]~q ;
wire \mem~12_combout ;
wire \mem[1][110]~q ;
wire \mem~13_combout ;
wire \mem[1][111]~q ;
wire \mem~14_combout ;
wire \mem[1][112]~q ;
wire \mem~15_combout ;
wire \mem[1][113]~q ;
wire \mem~16_combout ;
wire \mem[1][114]~q ;
wire \mem~17_combout ;
wire \mem[1][115]~q ;
wire \mem~18_combout ;
wire \mem[1][116]~q ;
wire \mem~19_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][129] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_129_0),
	.prn(vcc));
defparam \mem[0][129] .is_wysiwyg = "true";
defparam \mem[0][129] .power_up = "low";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][68] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_68_0),
	.prn(vcc));
defparam \mem[0][68] .is_wysiwyg = "true";
defparam \mem[0][68] .power_up = "low";

dffeas \mem[0][66] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_66_0),
	.prn(vcc));
defparam \mem[0][66] .is_wysiwyg = "true";
defparam \mem[0][66] .power_up = "low";

dffeas \mem[0][130] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_130_0),
	.prn(vcc));
defparam \mem[0][130] .is_wysiwyg = "true";
defparam \mem[0][130] .power_up = "low";

dffeas \mem[0][78] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_78_0),
	.prn(vcc));
defparam \mem[0][78] .is_wysiwyg = "true";
defparam \mem[0][78] .power_up = "low";

dffeas \mem[0][77] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_77_0),
	.prn(vcc));
defparam \mem[0][77] .is_wysiwyg = "true";
defparam \mem[0][77] .power_up = "low";

dffeas \mem[0][76] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_76_0),
	.prn(vcc));
defparam \mem[0][76] .is_wysiwyg = "true";
defparam \mem[0][76] .power_up = "low";

dffeas \mem[0][75] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_75_0),
	.prn(vcc));
defparam \mem[0][75] .is_wysiwyg = "true";
defparam \mem[0][75] .power_up = "low";

dffeas \mem[0][74] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_74_0),
	.prn(vcc));
defparam \mem[0][74] .is_wysiwyg = "true";
defparam \mem[0][74] .power_up = "low";

dffeas \mem[0][105] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_105_0),
	.prn(vcc));
defparam \mem[0][105] .is_wysiwyg = "true";
defparam \mem[0][105] .power_up = "low";

dffeas \mem[0][106] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_106_0),
	.prn(vcc));
defparam \mem[0][106] .is_wysiwyg = "true";
defparam \mem[0][106] .power_up = "low";

dffeas \mem[0][107] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_107_0),
	.prn(vcc));
defparam \mem[0][107] .is_wysiwyg = "true";
defparam \mem[0][107] .power_up = "low";

dffeas \mem[0][108] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_108_0),
	.prn(vcc));
defparam \mem[0][108] .is_wysiwyg = "true";
defparam \mem[0][108] .power_up = "low";

dffeas \mem[0][109] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_109_0),
	.prn(vcc));
defparam \mem[0][109] .is_wysiwyg = "true";
defparam \mem[0][109] .power_up = "low";

dffeas \mem[0][110] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_110_0),
	.prn(vcc));
defparam \mem[0][110] .is_wysiwyg = "true";
defparam \mem[0][110] .power_up = "low";

dffeas \mem[0][111] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_111_0),
	.prn(vcc));
defparam \mem[0][111] .is_wysiwyg = "true";
defparam \mem[0][111] .power_up = "low";

dffeas \mem[0][112] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_112_0),
	.prn(vcc));
defparam \mem[0][112] .is_wysiwyg = "true";
defparam \mem[0][112] .power_up = "low";

dffeas \mem[0][113] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_113_0),
	.prn(vcc));
defparam \mem[0][113] .is_wysiwyg = "true";
defparam \mem[0][113] .power_up = "low";

dffeas \mem[0][114] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_114_0),
	.prn(vcc));
defparam \mem[0][114] .is_wysiwyg = "true";
defparam \mem[0][114] .power_up = "low";

dffeas \mem[0][115] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_115_0),
	.prn(vcc));
defparam \mem[0][115] .is_wysiwyg = "true";
defparam \mem[0][115] .power_up = "low";

dffeas \mem[0][116] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_116_0),
	.prn(vcc));
defparam \mem[0][116] .is_wysiwyg = "true";
defparam \mem[0][116] .power_up = "low";

cyclonev_lcell_comb \read~0 (
	.dataa(!comb),
	.datab(!WideOr01),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h1111111111111111;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \write~0 (
	.dataa(!mem_used_1),
	.datab(!WideOr0),
	.datac(!cp_ready),
	.datad(!rf_source_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'h008A008A008A008A;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!last_packet_beat),
	.datad(!read),
	.datae(!\write~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'h5505335355053353;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][129] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][129]~q ),
	.prn(vcc));
defparam \mem[1][129] .is_wysiwyg = "true";
defparam \mem[1][129] .power_up = "low";

cyclonev_lcell_comb \mem~20 (
	.dataa(!WideOr0),
	.datab(!out_valid_reg),
	.datac(!\mem[1][129]~q ),
	.datad(!in_data_reg_68),
	.datae(!mem_used_1),
	.dataf(!nxt_out_eop),
	.datag(!in_data_reg_69),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~20 .extended_lut = "on";
defparam \mem~20 .lut_mask = 64'h02020F0F02330F0F;
defparam \mem~20 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!mem_used_0),
	.datab(!rp_valid),
	.datac(!last_packet_beat),
	.datad(!read),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hAAEAAAEAAAEAAAEA;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!rp_valid),
	.datad(!last_packet_beat),
	.datae(!read),
	.dataf(!\write~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'h33331333FFFFFFFF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem[1][68] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][68]~q ),
	.prn(vcc));
defparam \mem[1][68] .is_wysiwyg = "true";
defparam \mem[1][68] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!mem_used_1),
	.datab(!in_data_reg_68),
	.datac(!\mem[1][68]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h2727272727272727;
defparam \mem~0 .shared_arith = "off";

dffeas \mem[1][69] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][69]~q ),
	.prn(vcc));
defparam \mem[1][69] .is_wysiwyg = "true";
defparam \mem[1][69] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!mem_used_1),
	.datab(!in_data_reg_69),
	.datac(!\mem[1][69]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h2727272727272727;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[1][130] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][130]~q ),
	.prn(vcc));
defparam \mem[1][130] .is_wysiwyg = "true";
defparam \mem[1][130] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!mem_used_1),
	.datab(!nxt_out_eop),
	.datac(!\mem[1][130]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h2727272727272727;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[1][78] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][78]~q ),
	.prn(vcc));
defparam \mem[1][78] .is_wysiwyg = "true";
defparam \mem[1][78] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_6),
	.datad(!\mem[1][78]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h0257025702570257;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][77] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][77]~q ),
	.prn(vcc));
defparam \mem[1][77] .is_wysiwyg = "true";
defparam \mem[1][77] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\mem[1][77]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h0257025702570257;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][76] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][76]~q ),
	.prn(vcc));
defparam \mem[1][76] .is_wysiwyg = "true";
defparam \mem[1][76] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!\mem[1][76]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h0257025702570257;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][75] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][75]~q ),
	.prn(vcc));
defparam \mem[1][75] .is_wysiwyg = "true";
defparam \mem[1][75] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\mem[1][75]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h0257025702570257;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[1][74] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][74]~q ),
	.prn(vcc));
defparam \mem[1][74] .is_wysiwyg = "true";
defparam \mem[1][74] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_byte_cnt_reg_2),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(!\mem[1][74]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h082A5D7F082A5D7F;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[1][105] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][105]~q ),
	.prn(vcc));
defparam \mem[1][105] .is_wysiwyg = "true";
defparam \mem[1][105] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][105]~q ),
	.datac(!in_data_reg_105),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~8 .shared_arith = "off";

dffeas \mem[1][106] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][106]~q ),
	.prn(vcc));
defparam \mem[1][106] .is_wysiwyg = "true";
defparam \mem[1][106] .power_up = "low";

cyclonev_lcell_comb \mem~9 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][106]~q ),
	.datac(!in_data_reg_106),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~9 .extended_lut = "off";
defparam \mem~9 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~9 .shared_arith = "off";

dffeas \mem[1][107] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][107]~q ),
	.prn(vcc));
defparam \mem[1][107] .is_wysiwyg = "true";
defparam \mem[1][107] .power_up = "low";

cyclonev_lcell_comb \mem~10 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][107]~q ),
	.datac(!in_data_reg_107),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~10 .extended_lut = "off";
defparam \mem~10 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~10 .shared_arith = "off";

dffeas \mem[1][108] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][108]~q ),
	.prn(vcc));
defparam \mem[1][108] .is_wysiwyg = "true";
defparam \mem[1][108] .power_up = "low";

cyclonev_lcell_comb \mem~11 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][108]~q ),
	.datac(!in_data_reg_108),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~11 .extended_lut = "off";
defparam \mem~11 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~11 .shared_arith = "off";

dffeas \mem[1][109] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][109]~q ),
	.prn(vcc));
defparam \mem[1][109] .is_wysiwyg = "true";
defparam \mem[1][109] .power_up = "low";

cyclonev_lcell_comb \mem~12 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][109]~q ),
	.datac(!in_data_reg_109),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~12 .extended_lut = "off";
defparam \mem~12 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~12 .shared_arith = "off";

dffeas \mem[1][110] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][110]~q ),
	.prn(vcc));
defparam \mem[1][110] .is_wysiwyg = "true";
defparam \mem[1][110] .power_up = "low";

cyclonev_lcell_comb \mem~13 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][110]~q ),
	.datac(!in_data_reg_110),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~13 .extended_lut = "off";
defparam \mem~13 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~13 .shared_arith = "off";

dffeas \mem[1][111] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][111]~q ),
	.prn(vcc));
defparam \mem[1][111] .is_wysiwyg = "true";
defparam \mem[1][111] .power_up = "low";

cyclonev_lcell_comb \mem~14 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][111]~q ),
	.datac(!in_data_reg_111),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~14 .extended_lut = "off";
defparam \mem~14 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~14 .shared_arith = "off";

dffeas \mem[1][112] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][112]~q ),
	.prn(vcc));
defparam \mem[1][112] .is_wysiwyg = "true";
defparam \mem[1][112] .power_up = "low";

cyclonev_lcell_comb \mem~15 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][112]~q ),
	.datac(!in_data_reg_112),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~15 .extended_lut = "off";
defparam \mem~15 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~15 .shared_arith = "off";

dffeas \mem[1][113] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][113]~q ),
	.prn(vcc));
defparam \mem[1][113] .is_wysiwyg = "true";
defparam \mem[1][113] .power_up = "low";

cyclonev_lcell_comb \mem~16 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][113]~q ),
	.datac(!in_data_reg_113),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~16 .extended_lut = "off";
defparam \mem~16 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~16 .shared_arith = "off";

dffeas \mem[1][114] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][114]~q ),
	.prn(vcc));
defparam \mem[1][114] .is_wysiwyg = "true";
defparam \mem[1][114] .power_up = "low";

cyclonev_lcell_comb \mem~17 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][114]~q ),
	.datac(!in_data_reg_114),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~17 .extended_lut = "off";
defparam \mem~17 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~17 .shared_arith = "off";

dffeas \mem[1][115] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][115]~q ),
	.prn(vcc));
defparam \mem[1][115] .is_wysiwyg = "true";
defparam \mem[1][115] .power_up = "low";

cyclonev_lcell_comb \mem~18 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][115]~q ),
	.datac(!in_data_reg_115),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~18 .extended_lut = "off";
defparam \mem~18 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~18 .shared_arith = "off";

dffeas \mem[1][116] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][116]~q ),
	.prn(vcc));
defparam \mem[1][116] .is_wysiwyg = "true";
defparam \mem[1][116] .power_up = "low";

cyclonev_lcell_comb \mem~19 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][116]~q ),
	.datac(!in_data_reg_116),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~19 .extended_lut = "off";
defparam \mem~19 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~19 .shared_arith = "off";

endmodule

module spw_babasu_altera_avalon_sc_fifo_26 (
	h2f_RREADY_0,
	read_latency_shift_reg_0,
	mem_used_0,
	empty1,
	mem_0_0,
	av_readdata_pre_0,
	mem_1_0,
	av_readdata_pre_1,
	mem_2_0,
	av_readdata_pre_2,
	mem_3_0,
	av_readdata_pre_3,
	mem_4_0,
	av_readdata_pre_4,
	mem_5_0,
	av_readdata_pre_5,
	mem_6_0,
	av_readdata_pre_6,
	mem_7_0,
	av_readdata_pre_7,
	reset,
	clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_RREADY_0;
input 	read_latency_shift_reg_0;
output 	mem_used_0;
output 	empty1;
output 	mem_0_0;
input 	av_readdata_pre_0;
output 	mem_1_0;
input 	av_readdata_pre_1;
output 	mem_2_0;
input 	av_readdata_pre_2;
output 	mem_3_0;
input 	av_readdata_pre_3;
output 	mem_4_0;
input 	av_readdata_pre_4;
output 	mem_5_0;
input 	av_readdata_pre_5;
output 	mem_6_0;
input 	av_readdata_pre_6;
output 	mem_7_0;
input 	av_readdata_pre_7;
input 	reset;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[1]~1_combout ;
wire \mem_used[1]~q ;
wire \mem_used[0]~0_combout ;
wire \mem[1][0]~q ;
wire \mem~0_combout ;
wire \always0~0_combout ;
wire \mem[1][1]~q ;
wire \mem~1_combout ;
wire \mem[1][2]~q ;
wire \mem~2_combout ;
wire \mem[1][3]~q ;
wire \mem~3_combout ;
wire \mem[1][4]~q ;
wire \mem~4_combout ;
wire \mem[1][5]~q ;
wire \mem~5_combout ;
wire \mem[1][6]~q ;
wire \mem~6_combout ;
wire \mem[1][7]~q ;
wire \mem~7_combout ;


dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb empty(
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(empty1),
	.sumout(),
	.cout(),
	.shareout());
defparam empty.extended_lut = "off";
defparam empty.lut_mask = 64'h8888888888888888;
defparam empty.shared_arith = "off";

dffeas \mem[0][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_0_0),
	.prn(vcc));
defparam \mem[0][0] .is_wysiwyg = "true";
defparam \mem[0][0] .power_up = "low";

dffeas \mem[0][1] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_1_0),
	.prn(vcc));
defparam \mem[0][1] .is_wysiwyg = "true";
defparam \mem[0][1] .power_up = "low";

dffeas \mem[0][2] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_2_0),
	.prn(vcc));
defparam \mem[0][2] .is_wysiwyg = "true";
defparam \mem[0][2] .power_up = "low";

dffeas \mem[0][3] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_3_0),
	.prn(vcc));
defparam \mem[0][3] .is_wysiwyg = "true";
defparam \mem[0][3] .power_up = "low";

dffeas \mem[0][4] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_4_0),
	.prn(vcc));
defparam \mem[0][4] .is_wysiwyg = "true";
defparam \mem[0][4] .power_up = "low";

dffeas \mem[0][5] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_5_0),
	.prn(vcc));
defparam \mem[0][5] .is_wysiwyg = "true";
defparam \mem[0][5] .power_up = "low";

dffeas \mem[0][6] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_6_0),
	.prn(vcc));
defparam \mem[0][6] .is_wysiwyg = "true";
defparam \mem[0][6] .power_up = "low";

dffeas \mem[0][7] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_7_0),
	.prn(vcc));
defparam \mem[0][7] .is_wysiwyg = "true";
defparam \mem[0][7] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!h2f_RREADY_0),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem_used[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'h02EA02EA02EA02EA;
defparam \mem_used[1]~1 .shared_arith = "off";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[1]~q ),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~0 (
	.dataa(!h2f_RREADY_0),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem_used[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~0 .extended_lut = "off";
defparam \mem_used[0]~0 .lut_mask = 64'h2B1F2B1F2B1F2B1F;
defparam \mem_used[0]~0 .shared_arith = "off";

dffeas \mem[1][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][0]~q ),
	.prn(vcc));
defparam \mem[1][0] .is_wysiwyg = "true";
defparam \mem[1][0] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!av_readdata_pre_0),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h4747474747474747;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!h2f_RREADY_0),
	.datab(!mem_used_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \always0~0 .shared_arith = "off";

dffeas \mem[1][1] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][1]~q ),
	.prn(vcc));
defparam \mem[1][1] .is_wysiwyg = "true";
defparam \mem[1][1] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!av_readdata_pre_1),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h4747474747474747;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[1][2] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][2]~q ),
	.prn(vcc));
defparam \mem[1][2] .is_wysiwyg = "true";
defparam \mem[1][2] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!av_readdata_pre_2),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h4747474747474747;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[1][3] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][3]~q ),
	.prn(vcc));
defparam \mem[1][3] .is_wysiwyg = "true";
defparam \mem[1][3] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!av_readdata_pre_3),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h4747474747474747;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][4] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][4]~q ),
	.prn(vcc));
defparam \mem[1][4] .is_wysiwyg = "true";
defparam \mem[1][4] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!av_readdata_pre_4),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h4747474747474747;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][5] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][5]~q ),
	.prn(vcc));
defparam \mem[1][5] .is_wysiwyg = "true";
defparam \mem[1][5] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!av_readdata_pre_5),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][5]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h4747474747474747;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][6] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][6]~q ),
	.prn(vcc));
defparam \mem[1][6] .is_wysiwyg = "true";
defparam \mem[1][6] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!av_readdata_pre_6),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][6]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h4747474747474747;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[1][7] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][7]~q ),
	.prn(vcc));
defparam \mem[1][7] .is_wysiwyg = "true";
defparam \mem[1][7] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!av_readdata_pre_7),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h4747474747474747;
defparam \mem~7 .shared_arith = "off";

endmodule

module spw_babasu_altera_avalon_sc_fifo_27 (
	h2f_RREADY_0,
	waitrequest_reset_override,
	mem_used_1,
	in_data_reg_69,
	wait_latency_counter_1,
	wait_latency_counter_0,
	nxt_out_eop,
	out_valid_reg,
	stateST_UNCOMP_WR_SUBBURST,
	mem_130_0,
	empty,
	mem_66_0,
	mem_used_0,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	mem_105_0,
	mem_106_0,
	mem_107_0,
	mem_108_0,
	mem_109_0,
	mem_110_0,
	mem_111_0,
	mem_112_0,
	mem_113_0,
	mem_114_0,
	mem_115_0,
	mem_116_0,
	reset,
	last_packet_beat,
	write,
	write1,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_6,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_RREADY_0;
input 	waitrequest_reset_override;
output 	mem_used_1;
input 	in_data_reg_69;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	nxt_out_eop;
input 	out_valid_reg;
input 	stateST_UNCOMP_WR_SUBBURST;
output 	mem_130_0;
input 	empty;
output 	mem_66_0;
output 	mem_used_0;
output 	mem_78_0;
output 	mem_77_0;
output 	mem_76_0;
output 	mem_75_0;
output 	mem_74_0;
output 	mem_105_0;
output 	mem_106_0;
output 	mem_107_0;
output 	mem_108_0;
output 	mem_109_0;
output 	mem_110_0;
output 	mem_111_0;
output 	mem_112_0;
output 	mem_113_0;
output 	mem_114_0;
output 	mem_115_0;
output 	mem_116_0;
input 	reset;
input 	last_packet_beat;
output 	write;
output 	write1;
input 	out_byte_cnt_reg_2;
input 	out_uncomp_byte_cnt_reg_6;
input 	out_uncomp_byte_cnt_reg_5;
input 	out_uncomp_byte_cnt_reg_4;
input 	out_uncomp_byte_cnt_reg_3;
input 	out_uncomp_byte_cnt_reg_2;
input 	in_data_reg_105;
input 	in_data_reg_106;
input 	in_data_reg_107;
input 	in_data_reg_108;
input 	in_data_reg_109;
input 	in_data_reg_110;
input 	in_data_reg_111;
input 	in_data_reg_112;
input 	in_data_reg_113;
input 	in_data_reg_114;
input 	in_data_reg_115;
input 	in_data_reg_116;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read~0_combout ;
wire \mem_used[1]~0_combout ;
wire \mem[1][130]~q ;
wire \mem~0_combout ;
wire \always0~0_combout ;
wire \mem[1][69]~q ;
wire \mem~1_combout ;
wire \mem_used[0]~1_combout ;
wire \mem[1][78]~q ;
wire \mem~2_combout ;
wire \mem[1][77]~q ;
wire \mem~3_combout ;
wire \mem[1][76]~q ;
wire \mem~4_combout ;
wire \mem[1][75]~q ;
wire \mem~5_combout ;
wire \mem[1][74]~q ;
wire \mem~6_combout ;
wire \mem[1][105]~q ;
wire \mem~7_combout ;
wire \mem[1][106]~q ;
wire \mem~8_combout ;
wire \mem[1][107]~q ;
wire \mem~9_combout ;
wire \mem[1][108]~q ;
wire \mem~10_combout ;
wire \mem[1][109]~q ;
wire \mem~11_combout ;
wire \mem[1][110]~q ;
wire \mem~12_combout ;
wire \mem[1][111]~q ;
wire \mem~13_combout ;
wire \mem[1][112]~q ;
wire \mem~14_combout ;
wire \mem[1][113]~q ;
wire \mem~15_combout ;
wire \mem[1][114]~q ;
wire \mem~16_combout ;
wire \mem[1][115]~q ;
wire \mem~17_combout ;
wire \mem[1][116]~q ;
wire \mem~18_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][130] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_130_0),
	.prn(vcc));
defparam \mem[0][130] .is_wysiwyg = "true";
defparam \mem[0][130] .power_up = "low";

dffeas \mem[0][66] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_66_0),
	.prn(vcc));
defparam \mem[0][66] .is_wysiwyg = "true";
defparam \mem[0][66] .power_up = "low";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][78] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_78_0),
	.prn(vcc));
defparam \mem[0][78] .is_wysiwyg = "true";
defparam \mem[0][78] .power_up = "low";

dffeas \mem[0][77] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_77_0),
	.prn(vcc));
defparam \mem[0][77] .is_wysiwyg = "true";
defparam \mem[0][77] .power_up = "low";

dffeas \mem[0][76] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_76_0),
	.prn(vcc));
defparam \mem[0][76] .is_wysiwyg = "true";
defparam \mem[0][76] .power_up = "low";

dffeas \mem[0][75] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_75_0),
	.prn(vcc));
defparam \mem[0][75] .is_wysiwyg = "true";
defparam \mem[0][75] .power_up = "low";

dffeas \mem[0][74] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_74_0),
	.prn(vcc));
defparam \mem[0][74] .is_wysiwyg = "true";
defparam \mem[0][74] .power_up = "low";

dffeas \mem[0][105] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_105_0),
	.prn(vcc));
defparam \mem[0][105] .is_wysiwyg = "true";
defparam \mem[0][105] .power_up = "low";

dffeas \mem[0][106] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_106_0),
	.prn(vcc));
defparam \mem[0][106] .is_wysiwyg = "true";
defparam \mem[0][106] .power_up = "low";

dffeas \mem[0][107] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_107_0),
	.prn(vcc));
defparam \mem[0][107] .is_wysiwyg = "true";
defparam \mem[0][107] .power_up = "low";

dffeas \mem[0][108] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_108_0),
	.prn(vcc));
defparam \mem[0][108] .is_wysiwyg = "true";
defparam \mem[0][108] .power_up = "low";

dffeas \mem[0][109] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_109_0),
	.prn(vcc));
defparam \mem[0][109] .is_wysiwyg = "true";
defparam \mem[0][109] .power_up = "low";

dffeas \mem[0][110] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_110_0),
	.prn(vcc));
defparam \mem[0][110] .is_wysiwyg = "true";
defparam \mem[0][110] .power_up = "low";

dffeas \mem[0][111] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_111_0),
	.prn(vcc));
defparam \mem[0][111] .is_wysiwyg = "true";
defparam \mem[0][111] .power_up = "low";

dffeas \mem[0][112] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_112_0),
	.prn(vcc));
defparam \mem[0][112] .is_wysiwyg = "true";
defparam \mem[0][112] .power_up = "low";

dffeas \mem[0][113] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_113_0),
	.prn(vcc));
defparam \mem[0][113] .is_wysiwyg = "true";
defparam \mem[0][113] .power_up = "low";

dffeas \mem[0][114] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_114_0),
	.prn(vcc));
defparam \mem[0][114] .is_wysiwyg = "true";
defparam \mem[0][114] .power_up = "low";

dffeas \mem[0][115] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_115_0),
	.prn(vcc));
defparam \mem[0][115] .is_wysiwyg = "true";
defparam \mem[0][115] .power_up = "low";

dffeas \mem[0][116] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_116_0),
	.prn(vcc));
defparam \mem[0][116] .is_wysiwyg = "true";
defparam \mem[0][116] .power_up = "low";

cyclonev_lcell_comb \write~0 (
	.dataa(!waitrequest_reset_override),
	.datab(!in_data_reg_69),
	.datac(!mem_used_1),
	.datad(!out_valid_reg),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'h0010001000100010;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \write~1 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!write),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write1),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~1 .extended_lut = "off";
defparam \write~1 .lut_mask = 64'h0202020202020202;
defparam \write~1 .shared_arith = "off";

cyclonev_lcell_comb \read~0 (
	.dataa(!h2f_RREADY_0),
	.datab(!empty),
	.datac(!last_packet_beat),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h4040404040404040;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!\read~0_combout ),
	.datad(!write1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'h5431543154315431;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][130] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][130]~q ),
	.prn(vcc));
defparam \mem[1][130] .is_wysiwyg = "true";
defparam \mem[1][130] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!mem_used_1),
	.datab(!nxt_out_eop),
	.datac(!\mem[1][130]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h2727272727272727;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!mem_used_0),
	.datab(!\read~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \always0~0 .shared_arith = "off";

dffeas \mem[1][69] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][69]~q ),
	.prn(vcc));
defparam \mem[1][69] .is_wysiwyg = "true";
defparam \mem[1][69] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!in_data_reg_69),
	.datab(!mem_used_1),
	.datac(!\mem[1][69]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h4747474747474747;
defparam \mem~1 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!\read~0_combout ),
	.datad(!write1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'h31FF31FF31FF31FF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem[1][78] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][78]~q ),
	.prn(vcc));
defparam \mem[1][78] .is_wysiwyg = "true";
defparam \mem[1][78] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_6),
	.datad(!\mem[1][78]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h0257025702570257;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[1][77] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][77]~q ),
	.prn(vcc));
defparam \mem[1][77] .is_wysiwyg = "true";
defparam \mem[1][77] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\mem[1][77]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h0257025702570257;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][76] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][76]~q ),
	.prn(vcc));
defparam \mem[1][76] .is_wysiwyg = "true";
defparam \mem[1][76] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!\mem[1][76]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h0257025702570257;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][75] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][75]~q ),
	.prn(vcc));
defparam \mem[1][75] .is_wysiwyg = "true";
defparam \mem[1][75] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\mem[1][75]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h0257025702570257;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][74] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][74]~q ),
	.prn(vcc));
defparam \mem[1][74] .is_wysiwyg = "true";
defparam \mem[1][74] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_byte_cnt_reg_2),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(!\mem[1][74]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h082A5D7F082A5D7F;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[1][105] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][105]~q ),
	.prn(vcc));
defparam \mem[1][105] .is_wysiwyg = "true";
defparam \mem[1][105] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][105]~q ),
	.datac(!in_data_reg_105),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[1][106] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][106]~q ),
	.prn(vcc));
defparam \mem[1][106] .is_wysiwyg = "true";
defparam \mem[1][106] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][106]~q ),
	.datac(!in_data_reg_106),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~8 .shared_arith = "off";

dffeas \mem[1][107] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][107]~q ),
	.prn(vcc));
defparam \mem[1][107] .is_wysiwyg = "true";
defparam \mem[1][107] .power_up = "low";

cyclonev_lcell_comb \mem~9 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][107]~q ),
	.datac(!in_data_reg_107),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~9 .extended_lut = "off";
defparam \mem~9 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~9 .shared_arith = "off";

dffeas \mem[1][108] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][108]~q ),
	.prn(vcc));
defparam \mem[1][108] .is_wysiwyg = "true";
defparam \mem[1][108] .power_up = "low";

cyclonev_lcell_comb \mem~10 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][108]~q ),
	.datac(!in_data_reg_108),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~10 .extended_lut = "off";
defparam \mem~10 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~10 .shared_arith = "off";

dffeas \mem[1][109] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][109]~q ),
	.prn(vcc));
defparam \mem[1][109] .is_wysiwyg = "true";
defparam \mem[1][109] .power_up = "low";

cyclonev_lcell_comb \mem~11 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][109]~q ),
	.datac(!in_data_reg_109),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~11 .extended_lut = "off";
defparam \mem~11 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~11 .shared_arith = "off";

dffeas \mem[1][110] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][110]~q ),
	.prn(vcc));
defparam \mem[1][110] .is_wysiwyg = "true";
defparam \mem[1][110] .power_up = "low";

cyclonev_lcell_comb \mem~12 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][110]~q ),
	.datac(!in_data_reg_110),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~12 .extended_lut = "off";
defparam \mem~12 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~12 .shared_arith = "off";

dffeas \mem[1][111] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][111]~q ),
	.prn(vcc));
defparam \mem[1][111] .is_wysiwyg = "true";
defparam \mem[1][111] .power_up = "low";

cyclonev_lcell_comb \mem~13 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][111]~q ),
	.datac(!in_data_reg_111),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~13 .extended_lut = "off";
defparam \mem~13 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~13 .shared_arith = "off";

dffeas \mem[1][112] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][112]~q ),
	.prn(vcc));
defparam \mem[1][112] .is_wysiwyg = "true";
defparam \mem[1][112] .power_up = "low";

cyclonev_lcell_comb \mem~14 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][112]~q ),
	.datac(!in_data_reg_112),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~14 .extended_lut = "off";
defparam \mem~14 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~14 .shared_arith = "off";

dffeas \mem[1][113] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][113]~q ),
	.prn(vcc));
defparam \mem[1][113] .is_wysiwyg = "true";
defparam \mem[1][113] .power_up = "low";

cyclonev_lcell_comb \mem~15 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][113]~q ),
	.datac(!in_data_reg_113),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~15 .extended_lut = "off";
defparam \mem~15 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~15 .shared_arith = "off";

dffeas \mem[1][114] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][114]~q ),
	.prn(vcc));
defparam \mem[1][114] .is_wysiwyg = "true";
defparam \mem[1][114] .power_up = "low";

cyclonev_lcell_comb \mem~16 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][114]~q ),
	.datac(!in_data_reg_114),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~16 .extended_lut = "off";
defparam \mem~16 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~16 .shared_arith = "off";

dffeas \mem[1][115] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][115]~q ),
	.prn(vcc));
defparam \mem[1][115] .is_wysiwyg = "true";
defparam \mem[1][115] .power_up = "low";

cyclonev_lcell_comb \mem~17 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][115]~q ),
	.datac(!in_data_reg_115),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~17 .extended_lut = "off";
defparam \mem~17 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~17 .shared_arith = "off";

dffeas \mem[1][116] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][116]~q ),
	.prn(vcc));
defparam \mem[1][116] .is_wysiwyg = "true";
defparam \mem[1][116] .power_up = "low";

cyclonev_lcell_comb \mem~18 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][116]~q ),
	.datac(!in_data_reg_116),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~18 .extended_lut = "off";
defparam \mem~18 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~18 .shared_arith = "off";

endmodule

module spw_babasu_altera_avalon_sc_fifo_28 (
	read_latency_shift_reg_0,
	mem_used_0,
	mem_129_0,
	mem_used_01,
	av_readdata_pre_0,
	always4,
	mem_0_0,
	av_readdata_pre_1,
	mem_1_0,
	av_readdata_pre_2,
	mem_2_0,
	av_readdata_pre_3,
	mem_3_0,
	av_readdata_pre_4,
	mem_4_0,
	av_readdata_pre_5,
	mem_5_0,
	av_readdata_pre_6,
	mem_6_0,
	reset,
	WideOr0,
	clk)/* synthesis synthesis_greybox=0 */;
input 	read_latency_shift_reg_0;
output 	mem_used_0;
input 	mem_129_0;
input 	mem_used_01;
input 	av_readdata_pre_0;
output 	always4;
output 	mem_0_0;
input 	av_readdata_pre_1;
output 	mem_1_0;
input 	av_readdata_pre_2;
output 	mem_2_0;
input 	av_readdata_pre_3;
output 	mem_3_0;
input 	av_readdata_pre_4;
output 	mem_4_0;
input 	av_readdata_pre_5;
output 	mem_5_0;
input 	av_readdata_pre_6;
output 	mem_6_0;
input 	reset;
input 	WideOr0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~q ;
wire \mem_used[0]~0_combout ;
wire \mem[1][0]~q ;
wire \mem~0_combout ;
wire \always0~0_combout ;
wire \mem[1][1]~q ;
wire \mem~1_combout ;
wire \mem[1][2]~q ;
wire \mem~2_combout ;
wire \mem[1][3]~q ;
wire \mem~3_combout ;
wire \mem[1][4]~q ;
wire \mem~4_combout ;
wire \mem[1][5]~q ;
wire \mem~5_combout ;
wire \mem[1][6]~q ;
wire \mem~6_combout ;


dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \always4~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always4),
	.sumout(),
	.cout(),
	.shareout());
defparam \always4~0 .extended_lut = "off";
defparam \always4~0 .lut_mask = 64'h4444444444444444;
defparam \always4~0 .shared_arith = "off";

dffeas \mem[0][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_0_0),
	.prn(vcc));
defparam \mem[0][0] .is_wysiwyg = "true";
defparam \mem[0][0] .power_up = "low";

dffeas \mem[0][1] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_1_0),
	.prn(vcc));
defparam \mem[0][1] .is_wysiwyg = "true";
defparam \mem[0][1] .power_up = "low";

dffeas \mem[0][2] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_2_0),
	.prn(vcc));
defparam \mem[0][2] .is_wysiwyg = "true";
defparam \mem[0][2] .power_up = "low";

dffeas \mem[0][3] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_3_0),
	.prn(vcc));
defparam \mem[0][3] .is_wysiwyg = "true";
defparam \mem[0][3] .power_up = "low";

dffeas \mem[0][4] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_4_0),
	.prn(vcc));
defparam \mem[0][4] .is_wysiwyg = "true";
defparam \mem[0][4] .power_up = "low";

dffeas \mem[0][5] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_5_0),
	.prn(vcc));
defparam \mem[0][5] .is_wysiwyg = "true";
defparam \mem[0][5] .power_up = "low";

dffeas \mem[0][6] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_6_0),
	.prn(vcc));
defparam \mem[0][6] .is_wysiwyg = "true";
defparam \mem[0][6] .power_up = "low";

cyclonev_lcell_comb \read~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_129_0),
	.datad(!mem_used_01),
	.datae(!WideOr0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h0000777000007770;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!\mem_used[1]~q ),
	.datad(!\read~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'h1F001F001F001F00;
defparam \mem_used[1]~1 .shared_arith = "off";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[1]~q ),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!\mem_used[1]~q ),
	.datad(!\read~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~0 .extended_lut = "off";
defparam \mem_used[0]~0 .lut_mask = 64'h731F731F731F731F;
defparam \mem_used[0]~0 .shared_arith = "off";

dffeas \mem[1][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][0]~q ),
	.prn(vcc));
defparam \mem[1][0] .is_wysiwyg = "true";
defparam \mem[1][0] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!av_readdata_pre_0),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h4747474747474747;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!mem_used_0),
	.datab(!\read~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \always0~0 .shared_arith = "off";

dffeas \mem[1][1] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][1]~q ),
	.prn(vcc));
defparam \mem[1][1] .is_wysiwyg = "true";
defparam \mem[1][1] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!av_readdata_pre_1),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h4747474747474747;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[1][2] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][2]~q ),
	.prn(vcc));
defparam \mem[1][2] .is_wysiwyg = "true";
defparam \mem[1][2] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!av_readdata_pre_2),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h4747474747474747;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[1][3] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][3]~q ),
	.prn(vcc));
defparam \mem[1][3] .is_wysiwyg = "true";
defparam \mem[1][3] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!av_readdata_pre_3),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h4747474747474747;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][4] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][4]~q ),
	.prn(vcc));
defparam \mem[1][4] .is_wysiwyg = "true";
defparam \mem[1][4] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!av_readdata_pre_4),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h4747474747474747;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][5] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][5]~q ),
	.prn(vcc));
defparam \mem[1][5] .is_wysiwyg = "true";
defparam \mem[1][5] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!av_readdata_pre_5),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][5]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h4747474747474747;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][6] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][6]~q ),
	.prn(vcc));
defparam \mem[1][6] .is_wysiwyg = "true";
defparam \mem[1][6] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!av_readdata_pre_6),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][6]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h4747474747474747;
defparam \mem~6 .shared_arith = "off";

endmodule

module spw_babasu_altera_avalon_sc_fifo_29 (
	out_valid_reg,
	mem_used_1,
	WideOr0,
	in_data_reg_68,
	stateST_UNCOMP_WR_SUBBURST,
	mem_129_0,
	mem_used_0,
	mem_68_0,
	mem_66_0,
	comb,
	mem_130_0,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	mem_105_0,
	mem_106_0,
	mem_107_0,
	mem_108_0,
	mem_109_0,
	mem_110_0,
	mem_111_0,
	mem_112_0,
	mem_113_0,
	mem_114_0,
	mem_115_0,
	mem_116_0,
	reset,
	nxt_out_eop,
	last_packet_beat,
	WideOr01,
	read,
	cp_ready,
	in_data_reg_69,
	rf_source_valid,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_6,
	sink_ready,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	clk)/* synthesis synthesis_greybox=0 */;
input 	out_valid_reg;
output 	mem_used_1;
input 	WideOr0;
input 	in_data_reg_68;
input 	stateST_UNCOMP_WR_SUBBURST;
output 	mem_129_0;
output 	mem_used_0;
output 	mem_68_0;
output 	mem_66_0;
input 	comb;
output 	mem_130_0;
output 	mem_78_0;
output 	mem_77_0;
output 	mem_76_0;
output 	mem_75_0;
output 	mem_74_0;
output 	mem_105_0;
output 	mem_106_0;
output 	mem_107_0;
output 	mem_108_0;
output 	mem_109_0;
output 	mem_110_0;
output 	mem_111_0;
output 	mem_112_0;
output 	mem_113_0;
output 	mem_114_0;
output 	mem_115_0;
output 	mem_116_0;
input 	reset;
input 	nxt_out_eop;
input 	last_packet_beat;
input 	WideOr01;
output 	read;
input 	cp_ready;
input 	in_data_reg_69;
input 	rf_source_valid;
input 	out_byte_cnt_reg_2;
input 	out_uncomp_byte_cnt_reg_4;
input 	out_uncomp_byte_cnt_reg_3;
input 	out_uncomp_byte_cnt_reg_2;
input 	out_uncomp_byte_cnt_reg_5;
input 	out_uncomp_byte_cnt_reg_6;
input 	sink_ready;
input 	in_data_reg_105;
input 	in_data_reg_106;
input 	in_data_reg_107;
input 	in_data_reg_108;
input 	in_data_reg_109;
input 	in_data_reg_110;
input 	in_data_reg_111;
input 	in_data_reg_112;
input 	in_data_reg_113;
input 	in_data_reg_114;
input 	in_data_reg_115;
input 	in_data_reg_116;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \write~0_combout ;
wire \mem_used[1]~0_combout ;
wire \mem[1][129]~q ;
wire \mem~20_combout ;
wire \always0~0_combout ;
wire \mem_used[0]~1_combout ;
wire \mem[1][68]~q ;
wire \mem~0_combout ;
wire \mem[1][69]~q ;
wire \mem~1_combout ;
wire \mem[1][130]~q ;
wire \mem~2_combout ;
wire \mem[1][78]~q ;
wire \mem~3_combout ;
wire \mem[1][77]~q ;
wire \mem~4_combout ;
wire \mem[1][76]~q ;
wire \mem~5_combout ;
wire \mem[1][75]~q ;
wire \mem~6_combout ;
wire \mem[1][74]~q ;
wire \mem~7_combout ;
wire \mem[1][105]~q ;
wire \mem~8_combout ;
wire \mem[1][106]~q ;
wire \mem~9_combout ;
wire \mem[1][107]~q ;
wire \mem~10_combout ;
wire \mem[1][108]~q ;
wire \mem~11_combout ;
wire \mem[1][109]~q ;
wire \mem~12_combout ;
wire \mem[1][110]~q ;
wire \mem~13_combout ;
wire \mem[1][111]~q ;
wire \mem~14_combout ;
wire \mem[1][112]~q ;
wire \mem~15_combout ;
wire \mem[1][113]~q ;
wire \mem~16_combout ;
wire \mem[1][114]~q ;
wire \mem~17_combout ;
wire \mem[1][115]~q ;
wire \mem~18_combout ;
wire \mem[1][116]~q ;
wire \mem~19_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][129] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_129_0),
	.prn(vcc));
defparam \mem[0][129] .is_wysiwyg = "true";
defparam \mem[0][129] .power_up = "low";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][68] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_68_0),
	.prn(vcc));
defparam \mem[0][68] .is_wysiwyg = "true";
defparam \mem[0][68] .power_up = "low";

dffeas \mem[0][66] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_66_0),
	.prn(vcc));
defparam \mem[0][66] .is_wysiwyg = "true";
defparam \mem[0][66] .power_up = "low";

dffeas \mem[0][130] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_130_0),
	.prn(vcc));
defparam \mem[0][130] .is_wysiwyg = "true";
defparam \mem[0][130] .power_up = "low";

dffeas \mem[0][78] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_78_0),
	.prn(vcc));
defparam \mem[0][78] .is_wysiwyg = "true";
defparam \mem[0][78] .power_up = "low";

dffeas \mem[0][77] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_77_0),
	.prn(vcc));
defparam \mem[0][77] .is_wysiwyg = "true";
defparam \mem[0][77] .power_up = "low";

dffeas \mem[0][76] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_76_0),
	.prn(vcc));
defparam \mem[0][76] .is_wysiwyg = "true";
defparam \mem[0][76] .power_up = "low";

dffeas \mem[0][75] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_75_0),
	.prn(vcc));
defparam \mem[0][75] .is_wysiwyg = "true";
defparam \mem[0][75] .power_up = "low";

dffeas \mem[0][74] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_74_0),
	.prn(vcc));
defparam \mem[0][74] .is_wysiwyg = "true";
defparam \mem[0][74] .power_up = "low";

dffeas \mem[0][105] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_105_0),
	.prn(vcc));
defparam \mem[0][105] .is_wysiwyg = "true";
defparam \mem[0][105] .power_up = "low";

dffeas \mem[0][106] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_106_0),
	.prn(vcc));
defparam \mem[0][106] .is_wysiwyg = "true";
defparam \mem[0][106] .power_up = "low";

dffeas \mem[0][107] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_107_0),
	.prn(vcc));
defparam \mem[0][107] .is_wysiwyg = "true";
defparam \mem[0][107] .power_up = "low";

dffeas \mem[0][108] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_108_0),
	.prn(vcc));
defparam \mem[0][108] .is_wysiwyg = "true";
defparam \mem[0][108] .power_up = "low";

dffeas \mem[0][109] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_109_0),
	.prn(vcc));
defparam \mem[0][109] .is_wysiwyg = "true";
defparam \mem[0][109] .power_up = "low";

dffeas \mem[0][110] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_110_0),
	.prn(vcc));
defparam \mem[0][110] .is_wysiwyg = "true";
defparam \mem[0][110] .power_up = "low";

dffeas \mem[0][111] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_111_0),
	.prn(vcc));
defparam \mem[0][111] .is_wysiwyg = "true";
defparam \mem[0][111] .power_up = "low";

dffeas \mem[0][112] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_112_0),
	.prn(vcc));
defparam \mem[0][112] .is_wysiwyg = "true";
defparam \mem[0][112] .power_up = "low";

dffeas \mem[0][113] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_113_0),
	.prn(vcc));
defparam \mem[0][113] .is_wysiwyg = "true";
defparam \mem[0][113] .power_up = "low";

dffeas \mem[0][114] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_114_0),
	.prn(vcc));
defparam \mem[0][114] .is_wysiwyg = "true";
defparam \mem[0][114] .power_up = "low";

dffeas \mem[0][115] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_115_0),
	.prn(vcc));
defparam \mem[0][115] .is_wysiwyg = "true";
defparam \mem[0][115] .power_up = "low";

dffeas \mem[0][116] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_116_0),
	.prn(vcc));
defparam \mem[0][116] .is_wysiwyg = "true";
defparam \mem[0][116] .power_up = "low";

cyclonev_lcell_comb \read~0 (
	.dataa(!comb),
	.datab(!WideOr01),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h1111111111111111;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \write~0 (
	.dataa(!mem_used_1),
	.datab(!WideOr0),
	.datac(!cp_ready),
	.datad(!rf_source_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'h008A008A008A008A;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!last_packet_beat),
	.datad(!read),
	.datae(!\write~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'h5505335355053353;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][129] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][129]~q ),
	.prn(vcc));
defparam \mem[1][129] .is_wysiwyg = "true";
defparam \mem[1][129] .power_up = "low";

cyclonev_lcell_comb \mem~20 (
	.dataa(!WideOr0),
	.datab(!out_valid_reg),
	.datac(!\mem[1][129]~q ),
	.datad(!in_data_reg_68),
	.datae(!mem_used_1),
	.dataf(!nxt_out_eop),
	.datag(!in_data_reg_69),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~20 .extended_lut = "on";
defparam \mem~20 .lut_mask = 64'h02020F0F02330F0F;
defparam \mem~20 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!mem_used_0),
	.datab(!sink_ready),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!\write~0_combout ),
	.datad(!sink_ready),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'h3F1F3F1F3F1F3F1F;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem[1][68] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][68]~q ),
	.prn(vcc));
defparam \mem[1][68] .is_wysiwyg = "true";
defparam \mem[1][68] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!mem_used_1),
	.datab(!in_data_reg_68),
	.datac(!\mem[1][68]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h2727272727272727;
defparam \mem~0 .shared_arith = "off";

dffeas \mem[1][69] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][69]~q ),
	.prn(vcc));
defparam \mem[1][69] .is_wysiwyg = "true";
defparam \mem[1][69] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!mem_used_1),
	.datab(!in_data_reg_69),
	.datac(!\mem[1][69]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h2727272727272727;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[1][130] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][130]~q ),
	.prn(vcc));
defparam \mem[1][130] .is_wysiwyg = "true";
defparam \mem[1][130] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!mem_used_1),
	.datab(!nxt_out_eop),
	.datac(!\mem[1][130]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h2727272727272727;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[1][78] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][78]~q ),
	.prn(vcc));
defparam \mem[1][78] .is_wysiwyg = "true";
defparam \mem[1][78] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_6),
	.datad(!\mem[1][78]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h0257025702570257;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][77] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][77]~q ),
	.prn(vcc));
defparam \mem[1][77] .is_wysiwyg = "true";
defparam \mem[1][77] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\mem[1][77]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h0257025702570257;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][76] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][76]~q ),
	.prn(vcc));
defparam \mem[1][76] .is_wysiwyg = "true";
defparam \mem[1][76] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!\mem[1][76]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h0257025702570257;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][75] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][75]~q ),
	.prn(vcc));
defparam \mem[1][75] .is_wysiwyg = "true";
defparam \mem[1][75] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\mem[1][75]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h0257025702570257;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[1][74] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][74]~q ),
	.prn(vcc));
defparam \mem[1][74] .is_wysiwyg = "true";
defparam \mem[1][74] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_byte_cnt_reg_2),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(!\mem[1][74]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h082A5D7F082A5D7F;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[1][105] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][105]~q ),
	.prn(vcc));
defparam \mem[1][105] .is_wysiwyg = "true";
defparam \mem[1][105] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][105]~q ),
	.datac(!in_data_reg_105),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~8 .shared_arith = "off";

dffeas \mem[1][106] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][106]~q ),
	.prn(vcc));
defparam \mem[1][106] .is_wysiwyg = "true";
defparam \mem[1][106] .power_up = "low";

cyclonev_lcell_comb \mem~9 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][106]~q ),
	.datac(!in_data_reg_106),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~9 .extended_lut = "off";
defparam \mem~9 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~9 .shared_arith = "off";

dffeas \mem[1][107] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][107]~q ),
	.prn(vcc));
defparam \mem[1][107] .is_wysiwyg = "true";
defparam \mem[1][107] .power_up = "low";

cyclonev_lcell_comb \mem~10 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][107]~q ),
	.datac(!in_data_reg_107),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~10 .extended_lut = "off";
defparam \mem~10 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~10 .shared_arith = "off";

dffeas \mem[1][108] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][108]~q ),
	.prn(vcc));
defparam \mem[1][108] .is_wysiwyg = "true";
defparam \mem[1][108] .power_up = "low";

cyclonev_lcell_comb \mem~11 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][108]~q ),
	.datac(!in_data_reg_108),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~11 .extended_lut = "off";
defparam \mem~11 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~11 .shared_arith = "off";

dffeas \mem[1][109] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][109]~q ),
	.prn(vcc));
defparam \mem[1][109] .is_wysiwyg = "true";
defparam \mem[1][109] .power_up = "low";

cyclonev_lcell_comb \mem~12 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][109]~q ),
	.datac(!in_data_reg_109),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~12 .extended_lut = "off";
defparam \mem~12 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~12 .shared_arith = "off";

dffeas \mem[1][110] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][110]~q ),
	.prn(vcc));
defparam \mem[1][110] .is_wysiwyg = "true";
defparam \mem[1][110] .power_up = "low";

cyclonev_lcell_comb \mem~13 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][110]~q ),
	.datac(!in_data_reg_110),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~13 .extended_lut = "off";
defparam \mem~13 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~13 .shared_arith = "off";

dffeas \mem[1][111] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][111]~q ),
	.prn(vcc));
defparam \mem[1][111] .is_wysiwyg = "true";
defparam \mem[1][111] .power_up = "low";

cyclonev_lcell_comb \mem~14 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][111]~q ),
	.datac(!in_data_reg_111),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~14 .extended_lut = "off";
defparam \mem~14 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~14 .shared_arith = "off";

dffeas \mem[1][112] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][112]~q ),
	.prn(vcc));
defparam \mem[1][112] .is_wysiwyg = "true";
defparam \mem[1][112] .power_up = "low";

cyclonev_lcell_comb \mem~15 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][112]~q ),
	.datac(!in_data_reg_112),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~15 .extended_lut = "off";
defparam \mem~15 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~15 .shared_arith = "off";

dffeas \mem[1][113] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][113]~q ),
	.prn(vcc));
defparam \mem[1][113] .is_wysiwyg = "true";
defparam \mem[1][113] .power_up = "low";

cyclonev_lcell_comb \mem~16 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][113]~q ),
	.datac(!in_data_reg_113),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~16 .extended_lut = "off";
defparam \mem~16 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~16 .shared_arith = "off";

dffeas \mem[1][114] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][114]~q ),
	.prn(vcc));
defparam \mem[1][114] .is_wysiwyg = "true";
defparam \mem[1][114] .power_up = "low";

cyclonev_lcell_comb \mem~17 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][114]~q ),
	.datac(!in_data_reg_114),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~17 .extended_lut = "off";
defparam \mem~17 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~17 .shared_arith = "off";

dffeas \mem[1][115] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][115]~q ),
	.prn(vcc));
defparam \mem[1][115] .is_wysiwyg = "true";
defparam \mem[1][115] .power_up = "low";

cyclonev_lcell_comb \mem~18 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][115]~q ),
	.datac(!in_data_reg_115),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~18 .extended_lut = "off";
defparam \mem~18 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~18 .shared_arith = "off";

dffeas \mem[1][116] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][116]~q ),
	.prn(vcc));
defparam \mem[1][116] .is_wysiwyg = "true";
defparam \mem[1][116] .power_up = "low";

cyclonev_lcell_comb \mem~19 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][116]~q ),
	.datac(!in_data_reg_116),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~19 .extended_lut = "off";
defparam \mem~19 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~19 .shared_arith = "off";

endmodule

module spw_babasu_altera_avalon_sc_fifo_30 (
	h2f_RREADY_0,
	read_latency_shift_reg_0,
	mem_used_0,
	empty1,
	mem_0_0,
	av_readdata_pre_0,
	reset,
	clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_RREADY_0;
input 	read_latency_shift_reg_0;
output 	mem_used_0;
output 	empty1;
output 	mem_0_0;
input 	av_readdata_pre_0;
input 	reset;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[1]~1_combout ;
wire \mem_used[1]~q ;
wire \mem_used[0]~0_combout ;
wire \mem[1][0]~q ;
wire \mem~0_combout ;
wire \mem[0][0]~1_combout ;


dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb empty(
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(empty1),
	.sumout(),
	.cout(),
	.shareout());
defparam empty.extended_lut = "off";
defparam empty.lut_mask = 64'h8888888888888888;
defparam empty.shared_arith = "off";

dffeas \mem[0][0] (
	.clk(clk),
	.d(\mem[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_0_0),
	.prn(vcc));
defparam \mem[0][0] .is_wysiwyg = "true";
defparam \mem[0][0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!h2f_RREADY_0),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem_used[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'h02EA02EA02EA02EA;
defparam \mem_used[1]~1 .shared_arith = "off";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[1]~q ),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~0 (
	.dataa(!h2f_RREADY_0),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem_used[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~0 .extended_lut = "off";
defparam \mem_used[0]~0 .lut_mask = 64'h2B1F2B1F2B1F2B1F;
defparam \mem_used[0]~0 .shared_arith = "off";

dffeas \mem[1][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][0]~q ),
	.prn(vcc));
defparam \mem[1][0] .is_wysiwyg = "true";
defparam \mem[1][0] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!av_readdata_pre_0),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h4747474747474747;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \mem[0][0]~1 (
	.dataa(!h2f_RREADY_0),
	.datab(!mem_used_0),
	.datac(!mem_0_0),
	.datad(!\mem~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem[0][0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem[0][0]~1 .extended_lut = "off";
defparam \mem[0][0]~1 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \mem[0][0]~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_avalon_sc_fifo_31 (
	h2f_RREADY_0,
	waitrequest_reset_override,
	in_data_reg_69,
	mem_used_1,
	wait_latency_counter_1,
	wait_latency_counter_0,
	out_valid_reg,
	stateST_UNCOMP_WR_SUBBURST,
	empty,
	mem_66_0,
	mem_used_0,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	last_packet_beat,
	mem_130_0,
	mem_105_0,
	mem_106_0,
	mem_107_0,
	mem_108_0,
	mem_109_0,
	mem_110_0,
	mem_111_0,
	mem_112_0,
	mem_113_0,
	mem_114_0,
	mem_115_0,
	mem_116_0,
	reset,
	nxt_out_eop,
	out_byte_cnt_reg_2,
	write,
	write1,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_6,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_RREADY_0;
input 	waitrequest_reset_override;
input 	in_data_reg_69;
output 	mem_used_1;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	out_valid_reg;
input 	stateST_UNCOMP_WR_SUBBURST;
input 	empty;
output 	mem_66_0;
output 	mem_used_0;
output 	mem_78_0;
output 	mem_77_0;
output 	mem_76_0;
output 	mem_75_0;
output 	mem_74_0;
input 	last_packet_beat;
output 	mem_130_0;
output 	mem_105_0;
output 	mem_106_0;
output 	mem_107_0;
output 	mem_108_0;
output 	mem_109_0;
output 	mem_110_0;
output 	mem_111_0;
output 	mem_112_0;
output 	mem_113_0;
output 	mem_114_0;
output 	mem_115_0;
output 	mem_116_0;
input 	reset;
input 	nxt_out_eop;
input 	out_byte_cnt_reg_2;
output 	write;
output 	write1;
input 	out_uncomp_byte_cnt_reg_3;
input 	out_uncomp_byte_cnt_reg_2;
input 	out_uncomp_byte_cnt_reg_6;
input 	out_uncomp_byte_cnt_reg_5;
input 	out_uncomp_byte_cnt_reg_4;
input 	in_data_reg_105;
input 	in_data_reg_106;
input 	in_data_reg_107;
input 	in_data_reg_108;
input 	in_data_reg_109;
input 	in_data_reg_110;
input 	in_data_reg_111;
input 	in_data_reg_112;
input 	in_data_reg_113;
input 	in_data_reg_114;
input 	in_data_reg_115;
input 	in_data_reg_116;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read~0_combout ;
wire \mem_used[1]~0_combout ;
wire \mem[1][69]~q ;
wire \mem~0_combout ;
wire \always0~0_combout ;
wire \mem_used[0]~1_combout ;
wire \mem[1][78]~q ;
wire \mem~1_combout ;
wire \mem[1][77]~q ;
wire \mem~2_combout ;
wire \mem[1][76]~q ;
wire \mem~3_combout ;
wire \mem[1][75]~q ;
wire \mem~4_combout ;
wire \mem[1][74]~q ;
wire \mem~5_combout ;
wire \mem[1][130]~q ;
wire \mem~6_combout ;
wire \mem[1][105]~q ;
wire \mem~7_combout ;
wire \mem[1][106]~q ;
wire \mem~8_combout ;
wire \mem[1][107]~q ;
wire \mem~9_combout ;
wire \mem[1][108]~q ;
wire \mem~10_combout ;
wire \mem[1][109]~q ;
wire \mem~11_combout ;
wire \mem[1][110]~q ;
wire \mem~12_combout ;
wire \mem[1][111]~q ;
wire \mem~13_combout ;
wire \mem[1][112]~q ;
wire \mem~14_combout ;
wire \mem[1][113]~q ;
wire \mem~15_combout ;
wire \mem[1][114]~q ;
wire \mem~16_combout ;
wire \mem[1][115]~q ;
wire \mem~17_combout ;
wire \mem[1][116]~q ;
wire \mem~18_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][66] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_66_0),
	.prn(vcc));
defparam \mem[0][66] .is_wysiwyg = "true";
defparam \mem[0][66] .power_up = "low";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][78] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_78_0),
	.prn(vcc));
defparam \mem[0][78] .is_wysiwyg = "true";
defparam \mem[0][78] .power_up = "low";

dffeas \mem[0][77] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_77_0),
	.prn(vcc));
defparam \mem[0][77] .is_wysiwyg = "true";
defparam \mem[0][77] .power_up = "low";

dffeas \mem[0][76] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_76_0),
	.prn(vcc));
defparam \mem[0][76] .is_wysiwyg = "true";
defparam \mem[0][76] .power_up = "low";

dffeas \mem[0][75] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_75_0),
	.prn(vcc));
defparam \mem[0][75] .is_wysiwyg = "true";
defparam \mem[0][75] .power_up = "low";

dffeas \mem[0][74] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_74_0),
	.prn(vcc));
defparam \mem[0][74] .is_wysiwyg = "true";
defparam \mem[0][74] .power_up = "low";

dffeas \mem[0][130] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_130_0),
	.prn(vcc));
defparam \mem[0][130] .is_wysiwyg = "true";
defparam \mem[0][130] .power_up = "low";

dffeas \mem[0][105] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_105_0),
	.prn(vcc));
defparam \mem[0][105] .is_wysiwyg = "true";
defparam \mem[0][105] .power_up = "low";

dffeas \mem[0][106] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_106_0),
	.prn(vcc));
defparam \mem[0][106] .is_wysiwyg = "true";
defparam \mem[0][106] .power_up = "low";

dffeas \mem[0][107] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_107_0),
	.prn(vcc));
defparam \mem[0][107] .is_wysiwyg = "true";
defparam \mem[0][107] .power_up = "low";

dffeas \mem[0][108] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_108_0),
	.prn(vcc));
defparam \mem[0][108] .is_wysiwyg = "true";
defparam \mem[0][108] .power_up = "low";

dffeas \mem[0][109] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_109_0),
	.prn(vcc));
defparam \mem[0][109] .is_wysiwyg = "true";
defparam \mem[0][109] .power_up = "low";

dffeas \mem[0][110] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_110_0),
	.prn(vcc));
defparam \mem[0][110] .is_wysiwyg = "true";
defparam \mem[0][110] .power_up = "low";

dffeas \mem[0][111] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_111_0),
	.prn(vcc));
defparam \mem[0][111] .is_wysiwyg = "true";
defparam \mem[0][111] .power_up = "low";

dffeas \mem[0][112] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_112_0),
	.prn(vcc));
defparam \mem[0][112] .is_wysiwyg = "true";
defparam \mem[0][112] .power_up = "low";

dffeas \mem[0][113] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_113_0),
	.prn(vcc));
defparam \mem[0][113] .is_wysiwyg = "true";
defparam \mem[0][113] .power_up = "low";

dffeas \mem[0][114] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_114_0),
	.prn(vcc));
defparam \mem[0][114] .is_wysiwyg = "true";
defparam \mem[0][114] .power_up = "low";

dffeas \mem[0][115] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_115_0),
	.prn(vcc));
defparam \mem[0][115] .is_wysiwyg = "true";
defparam \mem[0][115] .power_up = "low";

dffeas \mem[0][116] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_116_0),
	.prn(vcc));
defparam \mem[0][116] .is_wysiwyg = "true";
defparam \mem[0][116] .power_up = "low";

cyclonev_lcell_comb \write~0 (
	.dataa(!waitrequest_reset_override),
	.datab(!in_data_reg_69),
	.datac(!mem_used_1),
	.datad(!out_valid_reg),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'h0010001000100010;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \write~1 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!write),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write1),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~1 .extended_lut = "off";
defparam \write~1 .lut_mask = 64'h0202020202020202;
defparam \write~1 .shared_arith = "off";

cyclonev_lcell_comb \read~0 (
	.dataa(!h2f_RREADY_0),
	.datab(!empty),
	.datac(!last_packet_beat),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h4040404040404040;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!\read~0_combout ),
	.datad(!write1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'h5431543154315431;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][69] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][69]~q ),
	.prn(vcc));
defparam \mem[1][69] .is_wysiwyg = "true";
defparam \mem[1][69] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!in_data_reg_69),
	.datab(!mem_used_1),
	.datac(!\mem[1][69]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h4747474747474747;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!mem_used_0),
	.datab(!\read~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!\read~0_combout ),
	.datad(!write1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'h31FF31FF31FF31FF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem[1][78] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][78]~q ),
	.prn(vcc));
defparam \mem[1][78] .is_wysiwyg = "true";
defparam \mem[1][78] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_6),
	.datad(!\mem[1][78]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h0257025702570257;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[1][77] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][77]~q ),
	.prn(vcc));
defparam \mem[1][77] .is_wysiwyg = "true";
defparam \mem[1][77] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\mem[1][77]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h0257025702570257;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[1][76] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][76]~q ),
	.prn(vcc));
defparam \mem[1][76] .is_wysiwyg = "true";
defparam \mem[1][76] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!\mem[1][76]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h0257025702570257;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][75] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][75]~q ),
	.prn(vcc));
defparam \mem[1][75] .is_wysiwyg = "true";
defparam \mem[1][75] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\mem[1][75]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h0257025702570257;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][74] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][74]~q ),
	.prn(vcc));
defparam \mem[1][74] .is_wysiwyg = "true";
defparam \mem[1][74] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_byte_cnt_reg_2),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(!\mem[1][74]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h082A5D7F082A5D7F;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][130] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][130]~q ),
	.prn(vcc));
defparam \mem[1][130] .is_wysiwyg = "true";
defparam \mem[1][130] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!mem_used_1),
	.datab(!nxt_out_eop),
	.datac(!\mem[1][130]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h2727272727272727;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[1][105] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][105]~q ),
	.prn(vcc));
defparam \mem[1][105] .is_wysiwyg = "true";
defparam \mem[1][105] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][105]~q ),
	.datac(!in_data_reg_105),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[1][106] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][106]~q ),
	.prn(vcc));
defparam \mem[1][106] .is_wysiwyg = "true";
defparam \mem[1][106] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][106]~q ),
	.datac(!in_data_reg_106),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~8 .shared_arith = "off";

dffeas \mem[1][107] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][107]~q ),
	.prn(vcc));
defparam \mem[1][107] .is_wysiwyg = "true";
defparam \mem[1][107] .power_up = "low";

cyclonev_lcell_comb \mem~9 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][107]~q ),
	.datac(!in_data_reg_107),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~9 .extended_lut = "off";
defparam \mem~9 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~9 .shared_arith = "off";

dffeas \mem[1][108] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][108]~q ),
	.prn(vcc));
defparam \mem[1][108] .is_wysiwyg = "true";
defparam \mem[1][108] .power_up = "low";

cyclonev_lcell_comb \mem~10 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][108]~q ),
	.datac(!in_data_reg_108),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~10 .extended_lut = "off";
defparam \mem~10 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~10 .shared_arith = "off";

dffeas \mem[1][109] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][109]~q ),
	.prn(vcc));
defparam \mem[1][109] .is_wysiwyg = "true";
defparam \mem[1][109] .power_up = "low";

cyclonev_lcell_comb \mem~11 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][109]~q ),
	.datac(!in_data_reg_109),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~11 .extended_lut = "off";
defparam \mem~11 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~11 .shared_arith = "off";

dffeas \mem[1][110] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][110]~q ),
	.prn(vcc));
defparam \mem[1][110] .is_wysiwyg = "true";
defparam \mem[1][110] .power_up = "low";

cyclonev_lcell_comb \mem~12 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][110]~q ),
	.datac(!in_data_reg_110),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~12 .extended_lut = "off";
defparam \mem~12 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~12 .shared_arith = "off";

dffeas \mem[1][111] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][111]~q ),
	.prn(vcc));
defparam \mem[1][111] .is_wysiwyg = "true";
defparam \mem[1][111] .power_up = "low";

cyclonev_lcell_comb \mem~13 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][111]~q ),
	.datac(!in_data_reg_111),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~13 .extended_lut = "off";
defparam \mem~13 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~13 .shared_arith = "off";

dffeas \mem[1][112] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][112]~q ),
	.prn(vcc));
defparam \mem[1][112] .is_wysiwyg = "true";
defparam \mem[1][112] .power_up = "low";

cyclonev_lcell_comb \mem~14 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][112]~q ),
	.datac(!in_data_reg_112),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~14 .extended_lut = "off";
defparam \mem~14 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~14 .shared_arith = "off";

dffeas \mem[1][113] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][113]~q ),
	.prn(vcc));
defparam \mem[1][113] .is_wysiwyg = "true";
defparam \mem[1][113] .power_up = "low";

cyclonev_lcell_comb \mem~15 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][113]~q ),
	.datac(!in_data_reg_113),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~15 .extended_lut = "off";
defparam \mem~15 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~15 .shared_arith = "off";

dffeas \mem[1][114] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][114]~q ),
	.prn(vcc));
defparam \mem[1][114] .is_wysiwyg = "true";
defparam \mem[1][114] .power_up = "low";

cyclonev_lcell_comb \mem~16 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][114]~q ),
	.datac(!in_data_reg_114),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~16 .extended_lut = "off";
defparam \mem~16 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~16 .shared_arith = "off";

dffeas \mem[1][115] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][115]~q ),
	.prn(vcc));
defparam \mem[1][115] .is_wysiwyg = "true";
defparam \mem[1][115] .power_up = "low";

cyclonev_lcell_comb \mem~17 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][115]~q ),
	.datac(!in_data_reg_115),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~17 .extended_lut = "off";
defparam \mem~17 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~17 .shared_arith = "off";

dffeas \mem[1][116] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][116]~q ),
	.prn(vcc));
defparam \mem[1][116] .is_wysiwyg = "true";
defparam \mem[1][116] .power_up = "low";

cyclonev_lcell_comb \mem~18 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][116]~q ),
	.datac(!in_data_reg_116),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~18 .extended_lut = "off";
defparam \mem~18 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~18 .shared_arith = "off";

endmodule

module spw_babasu_altera_avalon_sc_fifo_32 (
	read_latency_shift_reg_0,
	mem_used_0,
	mem_129_0,
	mem_used_01,
	av_readdata_pre_0,
	mem_0_0,
	reset,
	WideOr0,
	clk)/* synthesis synthesis_greybox=0 */;
input 	read_latency_shift_reg_0;
output 	mem_used_0;
input 	mem_129_0;
input 	mem_used_01;
input 	av_readdata_pre_0;
output 	mem_0_0;
input 	reset;
input 	WideOr0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~q ;
wire \mem_used[0]~0_combout ;
wire \mem[1][0]~q ;
wire \mem~0_combout ;
wire \mem[0][0]~1_combout ;


dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][0] (
	.clk(clk),
	.d(\mem[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_0_0),
	.prn(vcc));
defparam \mem[0][0] .is_wysiwyg = "true";
defparam \mem[0][0] .power_up = "low";

cyclonev_lcell_comb \read~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_129_0),
	.datad(!mem_used_01),
	.datae(!WideOr0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h0000777000007770;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!\mem_used[1]~q ),
	.datad(!\read~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'h1F001F001F001F00;
defparam \mem_used[1]~1 .shared_arith = "off";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[1]~q ),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!\mem_used[1]~q ),
	.datad(!\read~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~0 .extended_lut = "off";
defparam \mem_used[0]~0 .lut_mask = 64'h731F731F731F731F;
defparam \mem_used[0]~0 .shared_arith = "off";

dffeas \mem[1][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][0]~q ),
	.prn(vcc));
defparam \mem[1][0] .is_wysiwyg = "true";
defparam \mem[1][0] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!av_readdata_pre_0),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h4747474747474747;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \mem[0][0]~1 (
	.dataa(!mem_used_0),
	.datab(!mem_0_0),
	.datac(!\read~0_combout ),
	.datad(!\mem~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem[0][0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem[0][0]~1 .extended_lut = "off";
defparam \mem[0][0]~1 .lut_mask = 64'h10BF10BF10BF10BF;
defparam \mem[0][0]~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_avalon_sc_fifo_33 (
	out_valid_reg,
	mem_used_1,
	WideOr0,
	in_data_reg_68,
	stateST_UNCOMP_WR_SUBBURST,
	mem_129_0,
	mem_used_0,
	mem_68_0,
	mem_66_0,
	comb,
	mem_130_0,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	mem_105_0,
	mem_106_0,
	mem_107_0,
	mem_108_0,
	mem_109_0,
	mem_110_0,
	mem_111_0,
	mem_112_0,
	mem_113_0,
	mem_114_0,
	mem_115_0,
	mem_116_0,
	reset,
	nxt_out_eop,
	last_packet_beat,
	WideOr01,
	read,
	cp_ready,
	in_data_reg_69,
	rf_source_valid,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_6,
	sink_ready,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	clk)/* synthesis synthesis_greybox=0 */;
input 	out_valid_reg;
output 	mem_used_1;
input 	WideOr0;
input 	in_data_reg_68;
input 	stateST_UNCOMP_WR_SUBBURST;
output 	mem_129_0;
output 	mem_used_0;
output 	mem_68_0;
output 	mem_66_0;
input 	comb;
output 	mem_130_0;
output 	mem_78_0;
output 	mem_77_0;
output 	mem_76_0;
output 	mem_75_0;
output 	mem_74_0;
output 	mem_105_0;
output 	mem_106_0;
output 	mem_107_0;
output 	mem_108_0;
output 	mem_109_0;
output 	mem_110_0;
output 	mem_111_0;
output 	mem_112_0;
output 	mem_113_0;
output 	mem_114_0;
output 	mem_115_0;
output 	mem_116_0;
input 	reset;
input 	nxt_out_eop;
input 	last_packet_beat;
input 	WideOr01;
output 	read;
input 	cp_ready;
input 	in_data_reg_69;
input 	rf_source_valid;
input 	out_byte_cnt_reg_2;
input 	out_uncomp_byte_cnt_reg_4;
input 	out_uncomp_byte_cnt_reg_3;
input 	out_uncomp_byte_cnt_reg_2;
input 	out_uncomp_byte_cnt_reg_5;
input 	out_uncomp_byte_cnt_reg_6;
input 	sink_ready;
input 	in_data_reg_105;
input 	in_data_reg_106;
input 	in_data_reg_107;
input 	in_data_reg_108;
input 	in_data_reg_109;
input 	in_data_reg_110;
input 	in_data_reg_111;
input 	in_data_reg_112;
input 	in_data_reg_113;
input 	in_data_reg_114;
input 	in_data_reg_115;
input 	in_data_reg_116;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \write~0_combout ;
wire \mem_used[1]~0_combout ;
wire \mem[1][129]~q ;
wire \mem~20_combout ;
wire \always0~0_combout ;
wire \mem_used[0]~1_combout ;
wire \mem[1][68]~q ;
wire \mem~0_combout ;
wire \mem[1][69]~q ;
wire \mem~1_combout ;
wire \mem[1][130]~q ;
wire \mem~2_combout ;
wire \mem[1][78]~q ;
wire \mem~3_combout ;
wire \mem[1][77]~q ;
wire \mem~4_combout ;
wire \mem[1][76]~q ;
wire \mem~5_combout ;
wire \mem[1][75]~q ;
wire \mem~6_combout ;
wire \mem[1][74]~q ;
wire \mem~7_combout ;
wire \mem[1][105]~q ;
wire \mem~8_combout ;
wire \mem[1][106]~q ;
wire \mem~9_combout ;
wire \mem[1][107]~q ;
wire \mem~10_combout ;
wire \mem[1][108]~q ;
wire \mem~11_combout ;
wire \mem[1][109]~q ;
wire \mem~12_combout ;
wire \mem[1][110]~q ;
wire \mem~13_combout ;
wire \mem[1][111]~q ;
wire \mem~14_combout ;
wire \mem[1][112]~q ;
wire \mem~15_combout ;
wire \mem[1][113]~q ;
wire \mem~16_combout ;
wire \mem[1][114]~q ;
wire \mem~17_combout ;
wire \mem[1][115]~q ;
wire \mem~18_combout ;
wire \mem[1][116]~q ;
wire \mem~19_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][129] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_129_0),
	.prn(vcc));
defparam \mem[0][129] .is_wysiwyg = "true";
defparam \mem[0][129] .power_up = "low";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][68] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_68_0),
	.prn(vcc));
defparam \mem[0][68] .is_wysiwyg = "true";
defparam \mem[0][68] .power_up = "low";

dffeas \mem[0][66] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_66_0),
	.prn(vcc));
defparam \mem[0][66] .is_wysiwyg = "true";
defparam \mem[0][66] .power_up = "low";

dffeas \mem[0][130] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_130_0),
	.prn(vcc));
defparam \mem[0][130] .is_wysiwyg = "true";
defparam \mem[0][130] .power_up = "low";

dffeas \mem[0][78] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_78_0),
	.prn(vcc));
defparam \mem[0][78] .is_wysiwyg = "true";
defparam \mem[0][78] .power_up = "low";

dffeas \mem[0][77] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_77_0),
	.prn(vcc));
defparam \mem[0][77] .is_wysiwyg = "true";
defparam \mem[0][77] .power_up = "low";

dffeas \mem[0][76] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_76_0),
	.prn(vcc));
defparam \mem[0][76] .is_wysiwyg = "true";
defparam \mem[0][76] .power_up = "low";

dffeas \mem[0][75] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_75_0),
	.prn(vcc));
defparam \mem[0][75] .is_wysiwyg = "true";
defparam \mem[0][75] .power_up = "low";

dffeas \mem[0][74] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_74_0),
	.prn(vcc));
defparam \mem[0][74] .is_wysiwyg = "true";
defparam \mem[0][74] .power_up = "low";

dffeas \mem[0][105] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_105_0),
	.prn(vcc));
defparam \mem[0][105] .is_wysiwyg = "true";
defparam \mem[0][105] .power_up = "low";

dffeas \mem[0][106] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_106_0),
	.prn(vcc));
defparam \mem[0][106] .is_wysiwyg = "true";
defparam \mem[0][106] .power_up = "low";

dffeas \mem[0][107] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_107_0),
	.prn(vcc));
defparam \mem[0][107] .is_wysiwyg = "true";
defparam \mem[0][107] .power_up = "low";

dffeas \mem[0][108] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_108_0),
	.prn(vcc));
defparam \mem[0][108] .is_wysiwyg = "true";
defparam \mem[0][108] .power_up = "low";

dffeas \mem[0][109] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_109_0),
	.prn(vcc));
defparam \mem[0][109] .is_wysiwyg = "true";
defparam \mem[0][109] .power_up = "low";

dffeas \mem[0][110] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_110_0),
	.prn(vcc));
defparam \mem[0][110] .is_wysiwyg = "true";
defparam \mem[0][110] .power_up = "low";

dffeas \mem[0][111] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_111_0),
	.prn(vcc));
defparam \mem[0][111] .is_wysiwyg = "true";
defparam \mem[0][111] .power_up = "low";

dffeas \mem[0][112] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_112_0),
	.prn(vcc));
defparam \mem[0][112] .is_wysiwyg = "true";
defparam \mem[0][112] .power_up = "low";

dffeas \mem[0][113] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_113_0),
	.prn(vcc));
defparam \mem[0][113] .is_wysiwyg = "true";
defparam \mem[0][113] .power_up = "low";

dffeas \mem[0][114] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_114_0),
	.prn(vcc));
defparam \mem[0][114] .is_wysiwyg = "true";
defparam \mem[0][114] .power_up = "low";

dffeas \mem[0][115] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_115_0),
	.prn(vcc));
defparam \mem[0][115] .is_wysiwyg = "true";
defparam \mem[0][115] .power_up = "low";

dffeas \mem[0][116] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_116_0),
	.prn(vcc));
defparam \mem[0][116] .is_wysiwyg = "true";
defparam \mem[0][116] .power_up = "low";

cyclonev_lcell_comb \read~0 (
	.dataa(!comb),
	.datab(!WideOr01),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h1111111111111111;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \write~0 (
	.dataa(!mem_used_1),
	.datab(!WideOr0),
	.datac(!cp_ready),
	.datad(!rf_source_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'h008A008A008A008A;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!last_packet_beat),
	.datad(!read),
	.datae(!\write~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'h5505335355053353;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][129] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][129]~q ),
	.prn(vcc));
defparam \mem[1][129] .is_wysiwyg = "true";
defparam \mem[1][129] .power_up = "low";

cyclonev_lcell_comb \mem~20 (
	.dataa(!WideOr0),
	.datab(!out_valid_reg),
	.datac(!\mem[1][129]~q ),
	.datad(!in_data_reg_68),
	.datae(!mem_used_1),
	.dataf(!nxt_out_eop),
	.datag(!in_data_reg_69),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~20 .extended_lut = "on";
defparam \mem~20 .lut_mask = 64'h02020F0F02330F0F;
defparam \mem~20 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!mem_used_0),
	.datab(!sink_ready),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!\write~0_combout ),
	.datad(!sink_ready),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'h3F1F3F1F3F1F3F1F;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem[1][68] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][68]~q ),
	.prn(vcc));
defparam \mem[1][68] .is_wysiwyg = "true";
defparam \mem[1][68] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!mem_used_1),
	.datab(!in_data_reg_68),
	.datac(!\mem[1][68]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h2727272727272727;
defparam \mem~0 .shared_arith = "off";

dffeas \mem[1][69] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][69]~q ),
	.prn(vcc));
defparam \mem[1][69] .is_wysiwyg = "true";
defparam \mem[1][69] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!mem_used_1),
	.datab(!in_data_reg_69),
	.datac(!\mem[1][69]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h2727272727272727;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[1][130] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][130]~q ),
	.prn(vcc));
defparam \mem[1][130] .is_wysiwyg = "true";
defparam \mem[1][130] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!mem_used_1),
	.datab(!nxt_out_eop),
	.datac(!\mem[1][130]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h2727272727272727;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[1][78] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][78]~q ),
	.prn(vcc));
defparam \mem[1][78] .is_wysiwyg = "true";
defparam \mem[1][78] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_6),
	.datad(!\mem[1][78]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h0257025702570257;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][77] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][77]~q ),
	.prn(vcc));
defparam \mem[1][77] .is_wysiwyg = "true";
defparam \mem[1][77] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\mem[1][77]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h0257025702570257;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][76] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][76]~q ),
	.prn(vcc));
defparam \mem[1][76] .is_wysiwyg = "true";
defparam \mem[1][76] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!\mem[1][76]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h0257025702570257;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][75] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][75]~q ),
	.prn(vcc));
defparam \mem[1][75] .is_wysiwyg = "true";
defparam \mem[1][75] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\mem[1][75]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h0257025702570257;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[1][74] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][74]~q ),
	.prn(vcc));
defparam \mem[1][74] .is_wysiwyg = "true";
defparam \mem[1][74] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_byte_cnt_reg_2),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(!\mem[1][74]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h082A5D7F082A5D7F;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[1][105] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][105]~q ),
	.prn(vcc));
defparam \mem[1][105] .is_wysiwyg = "true";
defparam \mem[1][105] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][105]~q ),
	.datac(!in_data_reg_105),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~8 .shared_arith = "off";

dffeas \mem[1][106] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][106]~q ),
	.prn(vcc));
defparam \mem[1][106] .is_wysiwyg = "true";
defparam \mem[1][106] .power_up = "low";

cyclonev_lcell_comb \mem~9 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][106]~q ),
	.datac(!in_data_reg_106),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~9 .extended_lut = "off";
defparam \mem~9 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~9 .shared_arith = "off";

dffeas \mem[1][107] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][107]~q ),
	.prn(vcc));
defparam \mem[1][107] .is_wysiwyg = "true";
defparam \mem[1][107] .power_up = "low";

cyclonev_lcell_comb \mem~10 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][107]~q ),
	.datac(!in_data_reg_107),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~10 .extended_lut = "off";
defparam \mem~10 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~10 .shared_arith = "off";

dffeas \mem[1][108] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][108]~q ),
	.prn(vcc));
defparam \mem[1][108] .is_wysiwyg = "true";
defparam \mem[1][108] .power_up = "low";

cyclonev_lcell_comb \mem~11 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][108]~q ),
	.datac(!in_data_reg_108),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~11 .extended_lut = "off";
defparam \mem~11 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~11 .shared_arith = "off";

dffeas \mem[1][109] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][109]~q ),
	.prn(vcc));
defparam \mem[1][109] .is_wysiwyg = "true";
defparam \mem[1][109] .power_up = "low";

cyclonev_lcell_comb \mem~12 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][109]~q ),
	.datac(!in_data_reg_109),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~12 .extended_lut = "off";
defparam \mem~12 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~12 .shared_arith = "off";

dffeas \mem[1][110] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][110]~q ),
	.prn(vcc));
defparam \mem[1][110] .is_wysiwyg = "true";
defparam \mem[1][110] .power_up = "low";

cyclonev_lcell_comb \mem~13 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][110]~q ),
	.datac(!in_data_reg_110),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~13 .extended_lut = "off";
defparam \mem~13 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~13 .shared_arith = "off";

dffeas \mem[1][111] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][111]~q ),
	.prn(vcc));
defparam \mem[1][111] .is_wysiwyg = "true";
defparam \mem[1][111] .power_up = "low";

cyclonev_lcell_comb \mem~14 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][111]~q ),
	.datac(!in_data_reg_111),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~14 .extended_lut = "off";
defparam \mem~14 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~14 .shared_arith = "off";

dffeas \mem[1][112] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][112]~q ),
	.prn(vcc));
defparam \mem[1][112] .is_wysiwyg = "true";
defparam \mem[1][112] .power_up = "low";

cyclonev_lcell_comb \mem~15 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][112]~q ),
	.datac(!in_data_reg_112),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~15 .extended_lut = "off";
defparam \mem~15 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~15 .shared_arith = "off";

dffeas \mem[1][113] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][113]~q ),
	.prn(vcc));
defparam \mem[1][113] .is_wysiwyg = "true";
defparam \mem[1][113] .power_up = "low";

cyclonev_lcell_comb \mem~16 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][113]~q ),
	.datac(!in_data_reg_113),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~16 .extended_lut = "off";
defparam \mem~16 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~16 .shared_arith = "off";

dffeas \mem[1][114] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][114]~q ),
	.prn(vcc));
defparam \mem[1][114] .is_wysiwyg = "true";
defparam \mem[1][114] .power_up = "low";

cyclonev_lcell_comb \mem~17 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][114]~q ),
	.datac(!in_data_reg_114),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~17 .extended_lut = "off";
defparam \mem~17 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~17 .shared_arith = "off";

dffeas \mem[1][115] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][115]~q ),
	.prn(vcc));
defparam \mem[1][115] .is_wysiwyg = "true";
defparam \mem[1][115] .power_up = "low";

cyclonev_lcell_comb \mem~18 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][115]~q ),
	.datac(!in_data_reg_115),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~18 .extended_lut = "off";
defparam \mem~18 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~18 .shared_arith = "off";

dffeas \mem[1][116] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][116]~q ),
	.prn(vcc));
defparam \mem[1][116] .is_wysiwyg = "true";
defparam \mem[1][116] .power_up = "low";

cyclonev_lcell_comb \mem~19 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][116]~q ),
	.datac(!in_data_reg_116),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~19 .extended_lut = "off";
defparam \mem~19 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~19 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_axi_master_ni (
	h2f_AWVALID_0,
	h2f_WLAST_0,
	h2f_WVALID_0,
	h2f_ARBURST_0,
	h2f_ARBURST_1,
	h2f_ARLEN_0,
	h2f_ARLEN_1,
	h2f_ARLEN_2,
	h2f_ARLEN_3,
	h2f_ARSIZE_0,
	h2f_ARSIZE_1,
	h2f_ARSIZE_2,
	h2f_AWADDR_0,
	h2f_AWADDR_1,
	h2f_AWADDR_2,
	h2f_AWADDR_3,
	h2f_AWADDR_4,
	h2f_AWADDR_5,
	h2f_AWADDR_6,
	h2f_AWADDR_7,
	h2f_AWADDR_8,
	h2f_AWBURST_0,
	h2f_AWBURST_1,
	h2f_AWLEN_0,
	h2f_AWLEN_1,
	h2f_AWLEN_2,
	h2f_AWLEN_3,
	h2f_AWSIZE_0,
	h2f_AWSIZE_1,
	h2f_AWSIZE_2,
	address_burst_8,
	address_burst_7,
	address_burst_6,
	Add5,
	Add51,
	Add52,
	write_addr_data_both_valid1,
	sop_enable1,
	out_data_8,
	address_burst_5,
	out_data_5,
	address_burst_4,
	out_data_4,
	out_data_7,
	out_data_6,
	nonposted_cmd_accepted,
	altera_reset_synchronizer_int_chain_out,
	Decoder1,
	Add2,
	Add21,
	Add22,
	Add23,
	burst_bytecount_5,
	write_cp_data_77,
	burst_bytecount_6,
	write_cp_data_78,
	burst_bytecount_3,
	write_cp_data_75,
	burst_bytecount_2,
	write_cp_data_74,
	burst_bytecount_4,
	write_cp_data_76,
	Selector3,
	Selector10,
	Selector101,
	base_address_3,
	Selector4,
	Add3,
	Add31,
	Selector11,
	Selector111,
	base_address_2,
	Selector5,
	Add32,
	Selector12,
	out_data_1,
	out_data_0,
	Selector6,
	Selector13,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_AWVALID_0;
input 	h2f_WLAST_0;
input 	h2f_WVALID_0;
input 	h2f_ARBURST_0;
input 	h2f_ARBURST_1;
input 	h2f_ARLEN_0;
input 	h2f_ARLEN_1;
input 	h2f_ARLEN_2;
input 	h2f_ARLEN_3;
input 	h2f_ARSIZE_0;
input 	h2f_ARSIZE_1;
input 	h2f_ARSIZE_2;
input 	h2f_AWADDR_0;
input 	h2f_AWADDR_1;
input 	h2f_AWADDR_2;
input 	h2f_AWADDR_3;
input 	h2f_AWADDR_4;
input 	h2f_AWADDR_5;
input 	h2f_AWADDR_6;
input 	h2f_AWADDR_7;
input 	h2f_AWADDR_8;
input 	h2f_AWBURST_0;
input 	h2f_AWBURST_1;
input 	h2f_AWLEN_0;
input 	h2f_AWLEN_1;
input 	h2f_AWLEN_2;
input 	h2f_AWLEN_3;
input 	h2f_AWSIZE_0;
input 	h2f_AWSIZE_1;
input 	h2f_AWSIZE_2;
output 	address_burst_8;
output 	address_burst_7;
output 	address_burst_6;
output 	Add5;
output 	Add51;
output 	Add52;
output 	write_addr_data_both_valid1;
output 	sop_enable1;
output 	out_data_8;
output 	address_burst_5;
output 	out_data_5;
output 	address_burst_4;
output 	out_data_4;
output 	out_data_7;
output 	out_data_6;
input 	nonposted_cmd_accepted;
input 	altera_reset_synchronizer_int_chain_out;
output 	Decoder1;
output 	Add2;
output 	Add21;
output 	Add22;
output 	Add23;
output 	burst_bytecount_5;
output 	write_cp_data_77;
output 	burst_bytecount_6;
output 	write_cp_data_78;
output 	burst_bytecount_3;
output 	write_cp_data_75;
output 	burst_bytecount_2;
output 	write_cp_data_74;
output 	burst_bytecount_4;
output 	write_cp_data_76;
output 	Selector3;
output 	Selector10;
output 	Selector101;
output 	base_address_3;
output 	Selector4;
output 	Add3;
output 	Add31;
output 	Selector11;
output 	Selector111;
output 	base_address_2;
output 	Selector5;
output 	Add32;
output 	Selector12;
output 	out_data_1;
output 	out_data_0;
output 	Selector6;
output 	Selector13;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \LessThan14~0_combout ;
wire \align_address_to_size|Selector26~0_combout ;
wire \align_address_to_size|Decoder0~4_combout ;
wire \align_address_to_size|Decoder0~5_combout ;
wire \align_address_to_size|Decoder0~6_combout ;
wire \align_address_to_size|Decoder0~7_combout ;
wire \Add5~6 ;
wire \Add5~10 ;
wire \Decoder1~1_combout ;
wire \Decoder1~2_combout ;
wire \Decoder1~3_combout ;
wire \Decoder1~4_combout ;
wire \Add5~14 ;
wire \sop_enable~0_combout ;
wire \Add7~0_combout ;
wire \Add0~0_combout ;
wire \Add7~1_combout ;
wire \Add7~2_combout ;
wire \Add7~3_combout ;
wire \Add4~14 ;
wire \Add4~10 ;
wire \Add4~6 ;
wire \Add4~1_sumout ;
wire \Add3~0_combout ;
wire \log2ceil~0_combout ;
wire \Add1~0_combout ;
wire \Add1~1_combout ;
wire \Selector4~0_combout ;
wire \Add4~5_sumout ;
wire \Add4~9_sumout ;
wire \Selector5~0_combout ;
wire \Add4~13_sumout ;
wire \Add5~13_sumout ;
wire \Selector13~0_combout ;


spw_babasu_altera_merlin_address_alignment align_address_to_size(
	.h2f_AWADDR_0(h2f_AWADDR_0),
	.h2f_AWADDR_1(h2f_AWADDR_1),
	.h2f_AWADDR_2(h2f_AWADDR_2),
	.h2f_AWADDR_3(h2f_AWADDR_3),
	.h2f_AWADDR_4(h2f_AWADDR_4),
	.h2f_AWADDR_5(h2f_AWADDR_5),
	.h2f_AWADDR_6(h2f_AWADDR_6),
	.h2f_AWADDR_7(h2f_AWADDR_7),
	.h2f_AWADDR_8(h2f_AWADDR_8),
	.h2f_AWBURST_0(h2f_AWBURST_0),
	.h2f_AWBURST_1(h2f_AWBURST_1),
	.h2f_AWLEN_3(h2f_AWLEN_3),
	.h2f_AWSIZE_0(h2f_AWSIZE_0),
	.h2f_AWSIZE_1(h2f_AWSIZE_1),
	.h2f_AWSIZE_2(h2f_AWSIZE_2),
	.address_burst_8(address_burst_8),
	.address_burst_7(address_burst_7),
	.address_burst_6(address_burst_6),
	.sop_enable(sop_enable1),
	.out_data_8(out_data_8),
	.address_burst_5(address_burst_5),
	.out_data_5(out_data_5),
	.address_burst_4(address_burst_4),
	.out_data_4(out_data_4),
	.out_data_7(out_data_7),
	.out_data_6(out_data_6),
	.nonposted_cmd_accepted(nonposted_cmd_accepted),
	.reset(altera_reset_synchronizer_int_chain_out),
	.log2ceil(\log2ceil~0_combout ),
	.Add1(\Add1~0_combout ),
	.Add11(\Add1~1_combout ),
	.LessThan14(\LessThan14~0_combout ),
	.Selector26(\align_address_to_size|Selector26~0_combout ),
	.base_address_3(base_address_3),
	.Selector4(\Selector4~0_combout ),
	.base_address_2(base_address_2),
	.Decoder0(\align_address_to_size|Decoder0~4_combout ),
	.Decoder01(\align_address_to_size|Decoder0~5_combout ),
	.Decoder02(\align_address_to_size|Decoder0~6_combout ),
	.Selector5(\Selector5~0_combout ),
	.out_data_1(out_data_1),
	.Decoder03(\align_address_to_size|Decoder0~7_combout ),
	.out_data_0(out_data_0),
	.clk(clk_clk));

cyclonev_lcell_comb \LessThan14~0 (
	.dataa(!h2f_AWLEN_3),
	.datab(!h2f_AWSIZE_1),
	.datac(!h2f_AWSIZE_2),
	.datad(!\log2ceil~0_combout ),
	.datae(!\Add1~0_combout ),
	.dataf(!\Add1~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan14~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan14~0 .extended_lut = "off";
defparam \LessThan14~0 .lut_mask = 64'hE8A0A080A0808000;
defparam \LessThan14~0 .shared_arith = "off";

cyclonev_lcell_comb \Add5~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder1~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add5~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add5),
	.cout(),
	.shareout());
defparam \Add5~1 .extended_lut = "off";
defparam \Add5~1 .lut_mask = 64'h00000000000000FF;
defparam \Add5~1 .shared_arith = "off";

cyclonev_lcell_comb \Add5~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder1~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add5~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add51),
	.cout(\Add5~6 ),
	.shareout());
defparam \Add5~5 .extended_lut = "off";
defparam \Add5~5 .lut_mask = 64'h00000000000000FF;
defparam \Add5~5 .shared_arith = "off";

cyclonev_lcell_comb \Add5~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder1~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add5~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add52),
	.cout(\Add5~10 ),
	.shareout());
defparam \Add5~9 .extended_lut = "off";
defparam \Add5~9 .lut_mask = 64'h00000000000000FF;
defparam \Add5~9 .shared_arith = "off";

cyclonev_lcell_comb write_addr_data_both_valid(
	.dataa(!h2f_AWVALID_0),
	.datab(!h2f_WVALID_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_addr_data_both_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam write_addr_data_both_valid.extended_lut = "off";
defparam write_addr_data_both_valid.lut_mask = 64'h1111111111111111;
defparam write_addr_data_both_valid.shared_arith = "off";

dffeas sop_enable(
	.clk(clk_clk),
	.d(\sop_enable~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(nonposted_cmd_accepted),
	.q(sop_enable1),
	.prn(vcc));
defparam sop_enable.is_wysiwyg = "true";
defparam sop_enable.power_up = "low";

cyclonev_lcell_comb \Decoder1~0 (
	.dataa(!h2f_ARSIZE_1),
	.datab(!h2f_ARSIZE_2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Decoder1),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder1~0 .extended_lut = "off";
defparam \Decoder1~0 .lut_mask = 64'h8888888888888888;
defparam \Decoder1~0 .shared_arith = "off";

cyclonev_lcell_comb \Add2~0 (
	.dataa(!h2f_ARLEN_0),
	.datab(!h2f_ARLEN_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Add2),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add2~0 .extended_lut = "off";
defparam \Add2~0 .lut_mask = 64'h6666666666666666;
defparam \Add2~0 .shared_arith = "off";

cyclonev_lcell_comb \Add2~1 (
	.dataa(!h2f_ARLEN_0),
	.datab(!h2f_ARLEN_1),
	.datac(!h2f_ARLEN_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Add21),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add2~1 .extended_lut = "off";
defparam \Add2~1 .lut_mask = 64'h1E1E1E1E1E1E1E1E;
defparam \Add2~1 .shared_arith = "off";

cyclonev_lcell_comb \Add2~2 (
	.dataa(!h2f_ARLEN_0),
	.datab(!h2f_ARLEN_1),
	.datac(!h2f_ARLEN_2),
	.datad(!h2f_ARLEN_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Add22),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add2~2 .extended_lut = "off";
defparam \Add2~2 .lut_mask = 64'h01FE01FE01FE01FE;
defparam \Add2~2 .shared_arith = "off";

cyclonev_lcell_comb \Add2~3 (
	.dataa(!h2f_ARLEN_0),
	.datab(!h2f_ARLEN_1),
	.datac(!h2f_ARLEN_2),
	.datad(!h2f_ARLEN_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Add23),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add2~3 .extended_lut = "off";
defparam \Add2~3 .lut_mask = 64'h0001000100010001;
defparam \Add2~3 .shared_arith = "off";

dffeas \burst_bytecount[5] (
	.clk(clk_clk),
	.d(\Add7~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(nonposted_cmd_accepted),
	.q(burst_bytecount_5),
	.prn(vcc));
defparam \burst_bytecount[5] .is_wysiwyg = "true";
defparam \burst_bytecount[5] .power_up = "low";

cyclonev_lcell_comb \write_cp_data[77]~0 (
	.dataa(!h2f_AWLEN_3),
	.datab(!sop_enable1),
	.datac(!burst_bytecount_5),
	.datad(!\Add0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_cp_data_77),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_cp_data[77]~0 .extended_lut = "off";
defparam \write_cp_data[77]~0 .lut_mask = 64'h478B478B478B478B;
defparam \write_cp_data[77]~0 .shared_arith = "off";

dffeas \burst_bytecount[6] (
	.clk(clk_clk),
	.d(\Add7~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(nonposted_cmd_accepted),
	.q(burst_bytecount_6),
	.prn(vcc));
defparam \burst_bytecount[6] .is_wysiwyg = "true";
defparam \burst_bytecount[6] .power_up = "low";

cyclonev_lcell_comb \write_cp_data[78]~1 (
	.dataa(!h2f_AWLEN_3),
	.datab(!sop_enable1),
	.datac(!\Add0~0_combout ),
	.datad(!burst_bytecount_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_cp_data_78),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_cp_data[78]~1 .extended_lut = "off";
defparam \write_cp_data[78]~1 .lut_mask = 64'h0437043704370437;
defparam \write_cp_data[78]~1 .shared_arith = "off";

dffeas \burst_bytecount[3] (
	.clk(clk_clk),
	.d(\Add7~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(nonposted_cmd_accepted),
	.q(burst_bytecount_3),
	.prn(vcc));
defparam \burst_bytecount[3] .is_wysiwyg = "true";
defparam \burst_bytecount[3] .power_up = "low";

cyclonev_lcell_comb \write_cp_data[75]~2 (
	.dataa(!h2f_AWLEN_0),
	.datab(!h2f_AWLEN_1),
	.datac(!sop_enable1),
	.datad(!burst_bytecount_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_cp_data_75),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_cp_data[75]~2 .extended_lut = "off";
defparam \write_cp_data[75]~2 .lut_mask = 64'h606F606F606F606F;
defparam \write_cp_data[75]~2 .shared_arith = "off";

dffeas \burst_bytecount[2] (
	.clk(clk_clk),
	.d(write_cp_data_74),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(nonposted_cmd_accepted),
	.q(burst_bytecount_2),
	.prn(vcc));
defparam \burst_bytecount[2] .is_wysiwyg = "true";
defparam \burst_bytecount[2] .power_up = "low";

cyclonev_lcell_comb \write_cp_data[74]~3 (
	.dataa(!h2f_AWLEN_0),
	.datab(!sop_enable1),
	.datac(!burst_bytecount_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_cp_data_74),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_cp_data[74]~3 .extended_lut = "off";
defparam \write_cp_data[74]~3 .lut_mask = 64'h7474747474747474;
defparam \write_cp_data[74]~3 .shared_arith = "off";

dffeas \burst_bytecount[4] (
	.clk(clk_clk),
	.d(\Add7~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(nonposted_cmd_accepted),
	.q(burst_bytecount_4),
	.prn(vcc));
defparam \burst_bytecount[4] .is_wysiwyg = "true";
defparam \burst_bytecount[4] .power_up = "low";

cyclonev_lcell_comb \write_cp_data[76]~4 (
	.dataa(!h2f_AWLEN_0),
	.datab(!h2f_AWLEN_1),
	.datac(!h2f_AWLEN_2),
	.datad(!sop_enable1),
	.datae(!burst_bytecount_4),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_cp_data_76),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_cp_data[76]~4 .extended_lut = "off";
defparam \write_cp_data[76]~4 .lut_mask = 64'h1E001EFF1E001EFF;
defparam \write_cp_data[76]~4 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~0 (
	.dataa(!h2f_AWBURST_0),
	.datab(!h2f_AWBURST_1),
	.datac(!\Add4~1_sumout ),
	.datad(!\align_address_to_size|Selector26~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector3),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'h7F5D7F5D7F5D7F5D;
defparam \Selector3~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector10~0 (
	.dataa(!h2f_ARLEN_3),
	.datab(!h2f_ARSIZE_2),
	.datac(!\Add3~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector10),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector10~0 .extended_lut = "off";
defparam \Selector10~0 .lut_mask = 64'h8080808080808080;
defparam \Selector10~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector10~1 (
	.dataa(!h2f_ARBURST_0),
	.datab(!h2f_ARBURST_1),
	.datac(!Add5),
	.datad(!Selector10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector101),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector10~1 .extended_lut = "off";
defparam \Selector10~1 .lut_mask = 64'h7F5D7F5D7F5D7F5D;
defparam \Selector10~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector4~1 (
	.dataa(!h2f_AWBURST_0),
	.datab(!h2f_AWBURST_1),
	.datac(!\Selector4~0_combout ),
	.datad(!\Add4~5_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector4),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector4~1 .extended_lut = "off";
defparam \Selector4~1 .lut_mask = 64'h75FD75FD75FD75FD;
defparam \Selector4~1 .shared_arith = "off";

cyclonev_lcell_comb \Add3~1 (
	.dataa(!h2f_ARLEN_3),
	.datab(!h2f_ARSIZE_2),
	.datac(!\Add3~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Add3),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add3~1 .extended_lut = "off";
defparam \Add3~1 .lut_mask = 64'h1717171717171717;
defparam \Add3~1 .shared_arith = "off";

cyclonev_lcell_comb \Add3~2 (
	.dataa(!h2f_ARLEN_3),
	.datab(!h2f_ARSIZE_2),
	.datac(!\Add3~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Add31),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add3~2 .extended_lut = "off";
defparam \Add3~2 .lut_mask = 64'h6969696969696969;
defparam \Add3~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector11~0 (
	.dataa(!h2f_ARLEN_0),
	.datab(!h2f_ARLEN_1),
	.datac(!h2f_ARLEN_2),
	.datad(!h2f_ARLEN_3),
	.datae(!h2f_ARSIZE_0),
	.dataf(!h2f_ARSIZE_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector11),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector11~0 .extended_lut = "off";
defparam \Selector11~0 .lut_mask = 64'h0F003000400080FF;
defparam \Selector11~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector11~1 (
	.dataa(!h2f_ARBURST_0),
	.datab(!h2f_ARBURST_1),
	.datac(!Add3),
	.datad(!Add31),
	.datae(!Add51),
	.dataf(!Selector11),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector111),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector11~1 .extended_lut = "off";
defparam \Selector11~1 .lut_mask = 64'h5777DFFF7777FFFF;
defparam \Selector11~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector5~1 (
	.dataa(!h2f_AWBURST_0),
	.datab(!h2f_AWBURST_1),
	.datac(!\Add4~9_sumout ),
	.datad(!\Selector5~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector5),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~1 .extended_lut = "off";
defparam \Selector5~1 .lut_mask = 64'h7F5D7F5D7F5D7F5D;
defparam \Selector5~1 .shared_arith = "off";

cyclonev_lcell_comb \Add3~3 (
	.dataa(!h2f_ARLEN_0),
	.datab(!h2f_ARLEN_1),
	.datac(!h2f_ARLEN_2),
	.datad(!h2f_ARLEN_3),
	.datae(!h2f_ARSIZE_0),
	.dataf(!h2f_ARSIZE_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Add32),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add3~3 .extended_lut = "off";
defparam \Add3~3 .lut_mask = 64'h3F007000C0FF8FFF;
defparam \Add3~3 .shared_arith = "off";

cyclonev_lcell_comb \Selector12~0 (
	.dataa(!h2f_ARBURST_0),
	.datab(!h2f_ARBURST_1),
	.datac(!Add3),
	.datad(!Add31),
	.datae(!Add32),
	.dataf(!Add52),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector12),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector12~0 .extended_lut = "off";
defparam \Selector12~0 .lut_mask = 64'h57777777DFFFFFFF;
defparam \Selector12~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector6~0 (
	.dataa(!h2f_AWBURST_0),
	.datab(!h2f_AWBURST_1),
	.datac(!\Add1~1_combout ),
	.datad(!\Add4~13_sumout ),
	.datae(!\Selector5~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector6),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector6~0 .extended_lut = "off";
defparam \Selector6~0 .lut_mask = 64'h77FF57DF77FF57DF;
defparam \Selector6~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector13~1 (
	.dataa(!h2f_ARBURST_0),
	.datab(!h2f_ARBURST_1),
	.datac(!\Decoder1~4_combout ),
	.datad(!\Add5~13_sumout ),
	.datae(!\Selector13~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector13),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector13~1 .extended_lut = "off";
defparam \Selector13~1 .lut_mask = 64'h77FF75FD77FF75FD;
defparam \Selector13~1 .shared_arith = "off";

cyclonev_lcell_comb \Decoder1~1 (
	.dataa(!h2f_ARSIZE_0),
	.datab(!h2f_ARSIZE_1),
	.datac(!h2f_ARSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder1~1 .extended_lut = "off";
defparam \Decoder1~1 .lut_mask = 64'h1010101010101010;
defparam \Decoder1~1 .shared_arith = "off";

cyclonev_lcell_comb \Decoder1~2 (
	.dataa(!h2f_ARSIZE_0),
	.datab(!h2f_ARSIZE_1),
	.datac(!h2f_ARSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder1~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder1~2 .extended_lut = "off";
defparam \Decoder1~2 .lut_mask = 64'h2020202020202020;
defparam \Decoder1~2 .shared_arith = "off";

cyclonev_lcell_comb \Decoder1~3 (
	.dataa(!h2f_ARSIZE_0),
	.datab(!h2f_ARSIZE_1),
	.datac(!h2f_ARSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder1~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder1~3 .extended_lut = "off";
defparam \Decoder1~3 .lut_mask = 64'h4040404040404040;
defparam \Decoder1~3 .shared_arith = "off";

cyclonev_lcell_comb \Decoder1~4 (
	.dataa(!h2f_ARSIZE_0),
	.datab(!h2f_ARSIZE_1),
	.datac(!h2f_ARSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder1~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder1~4 .extended_lut = "off";
defparam \Decoder1~4 .lut_mask = 64'h8080808080808080;
defparam \Decoder1~4 .shared_arith = "off";

cyclonev_lcell_comb \Add5~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder1~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add5~13_sumout ),
	.cout(\Add5~14 ),
	.shareout());
defparam \Add5~13 .extended_lut = "off";
defparam \Add5~13 .lut_mask = 64'h00000000000000FF;
defparam \Add5~13 .shared_arith = "off";

cyclonev_lcell_comb \sop_enable~0 (
	.dataa(!h2f_WLAST_0),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sop_enable~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sop_enable~0 .extended_lut = "off";
defparam \sop_enable~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \sop_enable~0 .shared_arith = "off";

cyclonev_lcell_comb \Add7~0 (
	.dataa(!write_cp_data_74),
	.datab(!write_cp_data_75),
	.datac(!write_cp_data_76),
	.datad(!write_cp_data_77),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add7~0 .extended_lut = "off";
defparam \Add7~0 .lut_mask = 64'h40BF40BF40BF40BF;
defparam \Add7~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!h2f_AWLEN_0),
	.datab(!h2f_AWLEN_1),
	.datac(!h2f_AWLEN_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h0101010101010101;
defparam \Add0~0 .shared_arith = "off";

cyclonev_lcell_comb \Add7~1 (
	.dataa(!write_cp_data_74),
	.datab(!write_cp_data_75),
	.datac(!write_cp_data_76),
	.datad(!write_cp_data_77),
	.datae(!write_cp_data_78),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add7~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add7~1 .extended_lut = "off";
defparam \Add7~1 .lut_mask = 64'h4000BFFF4000BFFF;
defparam \Add7~1 .shared_arith = "off";

cyclonev_lcell_comb \Add7~2 (
	.dataa(!write_cp_data_74),
	.datab(!write_cp_data_75),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add7~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add7~2 .extended_lut = "off";
defparam \Add7~2 .lut_mask = 64'h6666666666666666;
defparam \Add7~2 .shared_arith = "off";

cyclonev_lcell_comb \Add7~3 (
	.dataa(!write_cp_data_74),
	.datab(!write_cp_data_75),
	.datac(!write_cp_data_76),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add7~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add7~3 .extended_lut = "off";
defparam \Add7~3 .lut_mask = 64'h4B4B4B4B4B4B4B4B;
defparam \Add7~3 .shared_arith = "off";

cyclonev_lcell_comb \Add4~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\align_address_to_size|Decoder0~7_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~13_sumout ),
	.cout(\Add4~14 ),
	.shareout());
defparam \Add4~13 .extended_lut = "off";
defparam \Add4~13 .lut_mask = 64'h00000000000000FF;
defparam \Add4~13 .shared_arith = "off";

cyclonev_lcell_comb \Add4~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\align_address_to_size|Decoder0~6_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~9_sumout ),
	.cout(\Add4~10 ),
	.shareout());
defparam \Add4~9 .extended_lut = "off";
defparam \Add4~9 .lut_mask = 64'h00000000000000FF;
defparam \Add4~9 .shared_arith = "off";

cyclonev_lcell_comb \Add4~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\align_address_to_size|Decoder0~5_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~5_sumout ),
	.cout(\Add4~6 ),
	.shareout());
defparam \Add4~5 .extended_lut = "off";
defparam \Add4~5 .lut_mask = 64'h00000000000000FF;
defparam \Add4~5 .shared_arith = "off";

cyclonev_lcell_comb \Add4~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\align_address_to_size|Decoder0~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~1_sumout ),
	.cout(),
	.shareout());
defparam \Add4~1 .extended_lut = "off";
defparam \Add4~1 .lut_mask = 64'h00000000000000FF;
defparam \Add4~1 .shared_arith = "off";

cyclonev_lcell_comb \Add3~0 (
	.dataa(!h2f_ARLEN_0),
	.datab(!h2f_ARLEN_1),
	.datac(!h2f_ARLEN_2),
	.datad(!h2f_ARLEN_3),
	.datae(!h2f_ARSIZE_0),
	.dataf(!h2f_ARSIZE_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add3~0 .extended_lut = "off";
defparam \Add3~0 .lut_mask = 64'h00000F003F007F00;
defparam \Add3~0 .shared_arith = "off";

cyclonev_lcell_comb \log2ceil~0 (
	.dataa(!h2f_AWLEN_1),
	.datab(!h2f_AWLEN_2),
	.datac(!h2f_AWLEN_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\log2ceil~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \log2ceil~0 .extended_lut = "off";
defparam \log2ceil~0 .lut_mask = 64'h7070707070707070;
defparam \log2ceil~0 .shared_arith = "off";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!h2f_AWLEN_0),
	.datab(!h2f_AWLEN_1),
	.datac(!h2f_AWLEN_2),
	.datad(!h2f_AWLEN_3),
	.datae(!h2f_AWSIZE_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h00004F0000004F00;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!h2f_AWLEN_0),
	.datab(!h2f_AWLEN_1),
	.datac(!h2f_AWLEN_2),
	.datad(!h2f_AWLEN_3),
	.datae(!h2f_AWSIZE_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h4F00B0FF4F00B0FF;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector4~0 (
	.dataa(!h2f_AWLEN_3),
	.datab(!h2f_AWSIZE_1),
	.datac(!h2f_AWSIZE_2),
	.datad(!\log2ceil~0_combout ),
	.datae(!\Add1~0_combout ),
	.dataf(!\Add1~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector4~0 .extended_lut = "off";
defparam \Selector4~0 .lut_mask = 64'hA080800080000000;
defparam \Selector4~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector5~0 (
	.dataa(!h2f_AWLEN_3),
	.datab(!h2f_AWSIZE_1),
	.datac(!h2f_AWSIZE_2),
	.datad(!\log2ceil~0_combout ),
	.datae(!\Add1~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~0 .extended_lut = "off";
defparam \Selector5~0 .lut_mask = 64'h8000000080000000;
defparam \Selector5~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector13~0 (
	.dataa(!h2f_ARLEN_0),
	.datab(!h2f_ARLEN_1),
	.datac(!h2f_ARLEN_2),
	.datad(!h2f_ARLEN_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector13~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector13~0 .extended_lut = "off";
defparam \Selector13~0 .lut_mask = 64'h8000800080008000;
defparam \Selector13~0 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_address_alignment (
	h2f_AWADDR_0,
	h2f_AWADDR_1,
	h2f_AWADDR_2,
	h2f_AWADDR_3,
	h2f_AWADDR_4,
	h2f_AWADDR_5,
	h2f_AWADDR_6,
	h2f_AWADDR_7,
	h2f_AWADDR_8,
	h2f_AWBURST_0,
	h2f_AWBURST_1,
	h2f_AWLEN_3,
	h2f_AWSIZE_0,
	h2f_AWSIZE_1,
	h2f_AWSIZE_2,
	address_burst_8,
	address_burst_7,
	address_burst_6,
	sop_enable,
	out_data_8,
	address_burst_5,
	out_data_5,
	address_burst_4,
	out_data_4,
	out_data_7,
	out_data_6,
	nonposted_cmd_accepted,
	reset,
	log2ceil,
	Add1,
	Add11,
	LessThan14,
	Selector26,
	base_address_3,
	Selector4,
	base_address_2,
	Decoder0,
	Decoder01,
	Decoder02,
	Selector5,
	out_data_1,
	Decoder03,
	out_data_0,
	clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_AWADDR_0;
input 	h2f_AWADDR_1;
input 	h2f_AWADDR_2;
input 	h2f_AWADDR_3;
input 	h2f_AWADDR_4;
input 	h2f_AWADDR_5;
input 	h2f_AWADDR_6;
input 	h2f_AWADDR_7;
input 	h2f_AWADDR_8;
input 	h2f_AWBURST_0;
input 	h2f_AWBURST_1;
input 	h2f_AWLEN_3;
input 	h2f_AWSIZE_0;
input 	h2f_AWSIZE_1;
input 	h2f_AWSIZE_2;
output 	address_burst_8;
output 	address_burst_7;
output 	address_burst_6;
input 	sop_enable;
output 	out_data_8;
output 	address_burst_5;
output 	out_data_5;
output 	address_burst_4;
output 	out_data_4;
output 	out_data_7;
output 	out_data_6;
input 	nonposted_cmd_accepted;
input 	reset;
input 	log2ceil;
input 	Add1;
input 	Add11;
input 	LessThan14;
output 	Selector26;
output 	base_address_3;
input 	Selector4;
output 	base_address_2;
output 	Decoder0;
output 	Decoder01;
output 	Decoder02;
input 	Selector5;
output 	out_data_1;
output 	Decoder03;
output 	out_data_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Decoder0~2_combout ;
wire \Decoder0~3_combout ;
wire \Decoder0~0_combout ;
wire \Decoder0~1_combout ;
wire \Add0~33_sumout ;
wire \Add1~21_sumout ;
wire \Selector29~0_combout ;
wire \address_burst[0]~q ;
wire \Add1~22 ;
wire \Add1~17_sumout ;
wire \aligned_address_bits[1]~combout ;
wire \Add0~34 ;
wire \Add0~29_sumout ;
wire \Selector28~0_combout ;
wire \address_burst[1]~q ;
wire \Add1~18 ;
wire \Add1~13_sumout ;
wire \Add0~30 ;
wire \Add0~25_sumout ;
wire \Selector27~0_combout ;
wire \address_burst[2]~q ;
wire \Add1~14 ;
wire \Add1~9_sumout ;
wire \Add0~26 ;
wire \Add0~21_sumout ;
wire \Selector26~1_combout ;
wire \address_burst[3]~q ;
wire \Add0~22 ;
wire \Add0~10 ;
wire \Add0~6 ;
wire \Add0~18 ;
wire \Add0~14 ;
wire \Add0~1_sumout ;
wire \Add0~13_sumout ;
wire \Add0~17_sumout ;
wire \Add1~10 ;
wire \Add1~6 ;
wire \Add1~1_sumout ;
wire \Selector24~0_combout ;
wire \Add0~5_sumout ;
wire \Selector24~1_combout ;
wire \Add1~5_sumout ;
wire \Add0~9_sumout ;
wire \Selector25~0_combout ;


dffeas \address_burst[8] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(out_data_8),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_AWBURST_0),
	.ena(nonposted_cmd_accepted),
	.q(address_burst_8),
	.prn(vcc));
defparam \address_burst[8] .is_wysiwyg = "true";
defparam \address_burst[8] .power_up = "low";

dffeas \address_burst[7] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(out_data_7),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_AWBURST_0),
	.ena(nonposted_cmd_accepted),
	.q(address_burst_7),
	.prn(vcc));
defparam \address_burst[7] .is_wysiwyg = "true";
defparam \address_burst[7] .power_up = "low";

dffeas \address_burst[6] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(out_data_6),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_AWBURST_0),
	.ena(nonposted_cmd_accepted),
	.q(address_burst_6),
	.prn(vcc));
defparam \address_burst[6] .is_wysiwyg = "true";
defparam \address_burst[6] .power_up = "low";

cyclonev_lcell_comb \out_data[8]~0 (
	.dataa(!h2f_AWADDR_8),
	.datab(!sop_enable),
	.datac(!address_burst_8),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[8]~0 .extended_lut = "off";
defparam \out_data[8]~0 .lut_mask = 64'h4747474747474747;
defparam \out_data[8]~0 .shared_arith = "off";

dffeas \address_burst[5] (
	.clk(clk),
	.d(\Selector24~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(nonposted_cmd_accepted),
	.q(address_burst_5),
	.prn(vcc));
defparam \address_burst[5] .is_wysiwyg = "true";
defparam \address_burst[5] .power_up = "low";

cyclonev_lcell_comb \out_data[5]~1 (
	.dataa(!h2f_AWADDR_5),
	.datab(!sop_enable),
	.datac(!address_burst_5),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[5]~1 .extended_lut = "off";
defparam \out_data[5]~1 .lut_mask = 64'h4747474747474747;
defparam \out_data[5]~1 .shared_arith = "off";

dffeas \address_burst[4] (
	.clk(clk),
	.d(\Selector25~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(nonposted_cmd_accepted),
	.q(address_burst_4),
	.prn(vcc));
defparam \address_burst[4] .is_wysiwyg = "true";
defparam \address_burst[4] .power_up = "low";

cyclonev_lcell_comb \out_data[4]~2 (
	.dataa(!h2f_AWADDR_4),
	.datab(!sop_enable),
	.datac(!address_burst_4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[4]~2 .extended_lut = "off";
defparam \out_data[4]~2 .lut_mask = 64'h4747474747474747;
defparam \out_data[4]~2 .shared_arith = "off";

cyclonev_lcell_comb \out_data[7]~3 (
	.dataa(!h2f_AWADDR_7),
	.datab(!sop_enable),
	.datac(!address_burst_7),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_7),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[7]~3 .extended_lut = "off";
defparam \out_data[7]~3 .lut_mask = 64'h4747474747474747;
defparam \out_data[7]~3 .shared_arith = "off";

cyclonev_lcell_comb \out_data[6]~4 (
	.dataa(!h2f_AWADDR_6),
	.datab(!sop_enable),
	.datac(!address_burst_6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_6),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[6]~4 .extended_lut = "off";
defparam \out_data[6]~4 .lut_mask = 64'h4747474747474747;
defparam \out_data[6]~4 .shared_arith = "off";

cyclonev_lcell_comb \Selector26~0 (
	.dataa(!h2f_AWLEN_3),
	.datab(!h2f_AWSIZE_1),
	.datac(!h2f_AWSIZE_2),
	.datad(!log2ceil),
	.datae(!Add1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector26),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector26~0 .extended_lut = "off";
defparam \Selector26~0 .lut_mask = 64'hA0808000A0808000;
defparam \Selector26~0 .shared_arith = "off";

cyclonev_lcell_comb \base_address[3]~0 (
	.dataa(!h2f_AWADDR_3),
	.datab(!sop_enable),
	.datac(!\address_burst[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(base_address_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \base_address[3]~0 .extended_lut = "off";
defparam \base_address[3]~0 .lut_mask = 64'h4747474747474747;
defparam \base_address[3]~0 .shared_arith = "off";

cyclonev_lcell_comb \base_address[2]~1 (
	.dataa(!h2f_AWADDR_2),
	.datab(!sop_enable),
	.datac(!\address_burst[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(base_address_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \base_address[2]~1 .extended_lut = "off";
defparam \base_address[2]~1 .lut_mask = 64'h4747474747474747;
defparam \base_address[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~4 (
	.dataa(!h2f_AWSIZE_0),
	.datab(!h2f_AWSIZE_1),
	.datac(!h2f_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Decoder0),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~4 .extended_lut = "off";
defparam \Decoder0~4 .lut_mask = 64'h1010101010101010;
defparam \Decoder0~4 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~5 (
	.dataa(!h2f_AWSIZE_0),
	.datab(!h2f_AWSIZE_1),
	.datac(!h2f_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Decoder01),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~5 .extended_lut = "off";
defparam \Decoder0~5 .lut_mask = 64'h2020202020202020;
defparam \Decoder0~5 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~6 (
	.dataa(!h2f_AWSIZE_0),
	.datab(!h2f_AWSIZE_1),
	.datac(!h2f_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Decoder02),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~6 .extended_lut = "off";
defparam \Decoder0~6 .lut_mask = 64'h4040404040404040;
defparam \Decoder0~6 .shared_arith = "off";

cyclonev_lcell_comb \out_data[1]~5 (
	.dataa(!h2f_AWADDR_1),
	.datab(!sop_enable),
	.datac(!\address_burst[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[1]~5 .extended_lut = "off";
defparam \out_data[1]~5 .lut_mask = 64'h4747474747474747;
defparam \out_data[1]~5 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~7 (
	.dataa(!h2f_AWSIZE_0),
	.datab(!h2f_AWSIZE_1),
	.datac(!h2f_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Decoder03),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~7 .extended_lut = "off";
defparam \Decoder0~7 .lut_mask = 64'h8080808080808080;
defparam \Decoder0~7 .shared_arith = "off";

cyclonev_lcell_comb \out_data[0]~6 (
	.dataa(!h2f_AWADDR_0),
	.datab(!sop_enable),
	.datac(!\address_burst[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[0]~6 .extended_lut = "off";
defparam \out_data[0]~6 .lut_mask = 64'h4747474747474747;
defparam \out_data[0]~6 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~2 (
	.dataa(!h2f_AWSIZE_0),
	.datab(!h2f_AWSIZE_1),
	.datac(!h2f_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~2 .extended_lut = "off";
defparam \Decoder0~2 .lut_mask = 64'h0101010101010101;
defparam \Decoder0~2 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~3 (
	.dataa(!h2f_AWSIZE_0),
	.datab(!h2f_AWSIZE_1),
	.datac(!h2f_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~3 .extended_lut = "off";
defparam \Decoder0~3 .lut_mask = 64'h0202020202020202;
defparam \Decoder0~3 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~0 (
	.dataa(!h2f_AWSIZE_0),
	.datab(!h2f_AWSIZE_1),
	.datac(!h2f_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~0 .extended_lut = "off";
defparam \Decoder0~0 .lut_mask = 64'h0404040404040404;
defparam \Decoder0~0 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~1 (
	.dataa(!h2f_AWSIZE_0),
	.datab(!h2f_AWSIZE_1),
	.datac(!h2f_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~1 .extended_lut = "off";
defparam \Decoder0~1 .lut_mask = 64'h0808080808080808;
defparam \Decoder0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~33 (
	.dataa(!sop_enable),
	.datab(!\address_burst[0]~q ),
	.datac(!h2f_AWADDR_0),
	.datad(!Decoder03),
	.datae(gnd),
	.dataf(!Decoder03),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h0000EEE4000000FF;
defparam \Add0~33 .shared_arith = "off";

cyclonev_lcell_comb \Add1~21 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!\address_burst[0]~q ),
	.datad(!Decoder03),
	.datae(gnd),
	.dataf(!h2f_AWADDR_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~21_sumout ),
	.cout(\Add1~22 ),
	.shareout());
defparam \Add1~21 .extended_lut = "off";
defparam \Add1~21 .lut_mask = 64'h0000FA50000000FF;
defparam \Add1~21 .shared_arith = "off";

cyclonev_lcell_comb \Selector29~0 (
	.dataa(!Add11),
	.datab(!out_data_0),
	.datac(!\Add0~33_sumout ),
	.datad(!\Add1~21_sumout ),
	.datae(!h2f_AWBURST_0),
	.dataf(!h2f_AWBURST_1),
	.datag(!Selector5),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector29~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector29~0 .extended_lut = "on";
defparam \Selector29~0 .lut_mask = 64'h33330F0F02F70F0F;
defparam \Selector29~0 .shared_arith = "off";

dffeas \address_burst[0] (
	.clk(clk),
	.d(\Selector29~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(nonposted_cmd_accepted),
	.q(\address_burst[0]~q ),
	.prn(vcc));
defparam \address_burst[0] .is_wysiwyg = "true";
defparam \address_burst[0] .power_up = "low";

cyclonev_lcell_comb \Add1~17 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!\address_burst[1]~q ),
	.datad(!Decoder02),
	.datae(gnd),
	.dataf(!h2f_AWADDR_1),
	.datag(gnd),
	.cin(\Add1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~17_sumout ),
	.cout(\Add1~18 ),
	.shareout());
defparam \Add1~17 .extended_lut = "off";
defparam \Add1~17 .lut_mask = 64'h0000FA50000000FF;
defparam \Add1~17 .shared_arith = "off";

cyclonev_lcell_comb \aligned_address_bits[1] (
	.dataa(!h2f_AWADDR_1),
	.datab(!h2f_AWSIZE_1),
	.datac(!h2f_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\aligned_address_bits[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \aligned_address_bits[1] .extended_lut = "off";
defparam \aligned_address_bits[1] .lut_mask = 64'h4040404040404040;
defparam \aligned_address_bits[1] .shared_arith = "off";

cyclonev_lcell_comb \Add0~29 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!\address_burst[1]~q ),
	.datad(!Decoder02),
	.datae(gnd),
	.dataf(!\aligned_address_bits[1]~combout ),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h0000FA50000000FF;
defparam \Add0~29 .shared_arith = "off";

cyclonev_lcell_comb \Selector28~0 (
	.dataa(!h2f_AWBURST_0),
	.datab(!h2f_AWBURST_1),
	.datac(!\Add1~17_sumout ),
	.datad(!\Add0~29_sumout ),
	.datae(!Selector5),
	.dataf(!out_data_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector28~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector28~0 .extended_lut = "off";
defparam \Selector28~0 .lut_mask = 64'h025700558ADFAAFF;
defparam \Selector28~0 .shared_arith = "off";

dffeas \address_burst[1] (
	.clk(clk),
	.d(\Selector28~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(nonposted_cmd_accepted),
	.q(\address_burst[1]~q ),
	.prn(vcc));
defparam \address_burst[1] .is_wysiwyg = "true";
defparam \address_burst[1] .power_up = "low";

cyclonev_lcell_comb \Add1~13 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_AWADDR_2),
	.datad(!Decoder01),
	.datae(gnd),
	.dataf(!\address_burst[2]~q ),
	.datag(gnd),
	.cin(\Add1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~13_sumout ),
	.cout(\Add1~14 ),
	.shareout());
defparam \Add1~13 .extended_lut = "off";
defparam \Add1~13 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add1~13 .shared_arith = "off";

cyclonev_lcell_comb \Add0~25 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_AWADDR_2),
	.datad(!Decoder01),
	.datae(gnd),
	.dataf(!\address_burst[2]~q ),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add0~25 .shared_arith = "off";

cyclonev_lcell_comb \Selector27~0 (
	.dataa(!h2f_AWBURST_0),
	.datab(!h2f_AWBURST_1),
	.datac(!Selector4),
	.datad(!base_address_2),
	.datae(!\Add1~13_sumout ),
	.dataf(!\Add0~25_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector27~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector27~0 .extended_lut = "off";
defparam \Selector27~0 .lut_mask = 64'h008A20AA55DF75FF;
defparam \Selector27~0 .shared_arith = "off";

dffeas \address_burst[2] (
	.clk(clk),
	.d(\Selector27~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(nonposted_cmd_accepted),
	.q(\address_burst[2]~q ),
	.prn(vcc));
defparam \address_burst[2] .is_wysiwyg = "true";
defparam \address_burst[2] .power_up = "low";

cyclonev_lcell_comb \Add1~9 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_AWADDR_3),
	.datad(!Decoder0),
	.datae(gnd),
	.dataf(!\address_burst[3]~q ),
	.datag(gnd),
	.cin(\Add1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~9_sumout ),
	.cout(\Add1~10 ),
	.shareout());
defparam \Add1~9 .extended_lut = "off";
defparam \Add1~9 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add1~9 .shared_arith = "off";

cyclonev_lcell_comb \Add0~21 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_AWADDR_3),
	.datad(!Decoder0),
	.datae(gnd),
	.dataf(!\address_burst[3]~q ),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add0~21 .shared_arith = "off";

cyclonev_lcell_comb \Selector26~1 (
	.dataa(!h2f_AWBURST_0),
	.datab(!h2f_AWBURST_1),
	.datac(!Selector26),
	.datad(!base_address_3),
	.datae(!\Add1~9_sumout ),
	.dataf(!\Add0~21_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector26~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector26~1 .extended_lut = "off";
defparam \Selector26~1 .lut_mask = 64'h008A20AA55DF75FF;
defparam \Selector26~1 .shared_arith = "off";

dffeas \address_burst[3] (
	.clk(clk),
	.d(\Selector26~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(nonposted_cmd_accepted),
	.q(\address_burst[3]~q ),
	.prn(vcc));
defparam \address_burst[3] .is_wysiwyg = "true";
defparam \address_burst[3] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_AWADDR_4),
	.datad(!\Decoder0~1_combout ),
	.datae(gnd),
	.dataf(!address_burst_4),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \Add0~5 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_AWADDR_5),
	.datad(!\Decoder0~0_combout ),
	.datae(gnd),
	.dataf(!address_burst_5),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~17 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_AWADDR_6),
	.datad(!\Decoder0~3_combout ),
	.datae(gnd),
	.dataf(!address_burst_6),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add0~17 .shared_arith = "off";

cyclonev_lcell_comb \Add0~13 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_AWADDR_7),
	.datad(!\Decoder0~2_combout ),
	.datae(gnd),
	.dataf(!address_burst_7),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_AWADDR_8),
	.datad(!address_burst_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FFFF00000A5F;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~5 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_AWADDR_4),
	.datad(!\Decoder0~1_combout ),
	.datae(gnd),
	.dataf(!address_burst_4),
	.datag(gnd),
	.cin(\Add1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~5_sumout ),
	.cout(\Add1~6 ),
	.shareout());
defparam \Add1~5 .extended_lut = "off";
defparam \Add1~5 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add1~5 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_AWADDR_5),
	.datad(!\Decoder0~0_combout ),
	.datae(gnd),
	.dataf(!address_burst_5),
	.datag(gnd),
	.cin(\Add1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~1_sumout ),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector24~0 (
	.dataa(!h2f_AWLEN_3),
	.datab(!h2f_AWSIZE_1),
	.datac(!h2f_AWSIZE_2),
	.datad(!log2ceil),
	.datae(!Add1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector24~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector24~0 .extended_lut = "off";
defparam \Selector24~0 .lut_mask = 64'hE8A0A080E8A0A080;
defparam \Selector24~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector24~1 (
	.dataa(!h2f_AWBURST_0),
	.datab(!h2f_AWBURST_1),
	.datac(!out_data_5),
	.datad(!\Add1~1_sumout ),
	.datae(!\Selector24~0_combout ),
	.dataf(!\Add0~5_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector24~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector24~1 .extended_lut = "off";
defparam \Selector24~1 .lut_mask = 64'h082A0A0A5D7F5F5F;
defparam \Selector24~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector25~0 (
	.dataa(!h2f_AWBURST_0),
	.datab(!h2f_AWBURST_1),
	.datac(!out_data_4),
	.datad(!\Add1~5_sumout ),
	.datae(!LessThan14),
	.dataf(!\Add0~9_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector25~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector25~0 .extended_lut = "off";
defparam \Selector25~0 .lut_mask = 64'h082A0A0A5D7F5F5F;
defparam \Selector25~0 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_burst_adapter (
	h2f_ARADDR_0,
	h2f_ARADDR_1,
	h2f_ARADDR_2,
	h2f_ARADDR_3,
	h2f_ARLEN_0,
	nxt_in_ready,
	in_ready_hold,
	stateST_COMP_TRANS,
	out_valid_reg,
	in_narrow_reg,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	in_data_reg_68,
	cp_ready,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready1,
	saved_grant_1,
	Equal16,
	saved_grant_0,
	in_data_reg_0,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	altera_reset_synchronizer_int_chain_out,
	Add2,
	Add21,
	Add22,
	Add23,
	write_cp_data_77,
	write_cp_data_78,
	write_cp_data_75,
	write_cp_data_74,
	write_cp_data_76,
	WideNor0,
	Equal14,
	nxt_out_eop,
	src2_valid,
	src_valid,
	cp_ready1,
	in_data_reg_69,
	src_data_87,
	src_data_88,
	src_valid1,
	src_data_35,
	src_data_34,
	src_data_33,
	src_data_32,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_6,
	src_payload_0,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	src_payload,
	Selector3,
	Selector10,
	src_data_82,
	base_address_3,
	Selector4,
	Selector11,
	src_data_81,
	base_address_2,
	src_data_105,
	src_data_106,
	src_data_107,
	src_data_108,
	src_data_109,
	src_data_110,
	src_data_111,
	src_data_112,
	src_data_113,
	src_data_114,
	src_data_115,
	src_data_116,
	src_data_86,
	Selector5,
	Selector12,
	src_data_80,
	out_data_1,
	out_data_0,
	Selector6,
	Selector13,
	src_data_79,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARADDR_0;
input 	h2f_ARADDR_1;
input 	h2f_ARADDR_2;
input 	h2f_ARADDR_3;
input 	h2f_ARLEN_0;
output 	nxt_in_ready;
output 	in_ready_hold;
output 	stateST_COMP_TRANS;
output 	out_valid_reg;
output 	in_narrow_reg;
output 	in_byteen_reg_3;
output 	in_byteen_reg_2;
output 	in_byteen_reg_1;
output 	in_byteen_reg_0;
output 	in_data_reg_68;
input 	cp_ready;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready1;
input 	saved_grant_1;
input 	Equal16;
input 	saved_grant_0;
output 	in_data_reg_0;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
input 	altera_reset_synchronizer_int_chain_out;
input 	Add2;
input 	Add21;
input 	Add22;
input 	Add23;
input 	write_cp_data_77;
input 	write_cp_data_78;
input 	write_cp_data_75;
input 	write_cp_data_74;
input 	write_cp_data_76;
input 	WideNor0;
input 	Equal14;
output 	nxt_out_eop;
input 	src2_valid;
input 	src_valid;
input 	cp_ready1;
output 	in_data_reg_69;
input 	src_data_87;
input 	src_data_88;
input 	src_valid1;
input 	src_data_35;
input 	src_data_34;
input 	src_data_33;
input 	src_data_32;
output 	out_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_6;
input 	src_payload_0;
output 	in_data_reg_105;
output 	in_data_reg_106;
output 	in_data_reg_107;
output 	in_data_reg_108;
output 	in_data_reg_109;
output 	in_data_reg_110;
output 	in_data_reg_111;
output 	in_data_reg_112;
output 	in_data_reg_113;
output 	in_data_reg_114;
output 	in_data_reg_115;
output 	in_data_reg_116;
input 	src_payload;
input 	Selector3;
input 	Selector10;
input 	src_data_82;
input 	base_address_3;
input 	Selector4;
input 	Selector11;
input 	src_data_81;
input 	base_address_2;
input 	src_data_105;
input 	src_data_106;
input 	src_data_107;
input 	src_data_108;
input 	src_data_109;
input 	src_data_110;
input 	src_data_111;
input 	src_data_112;
input 	src_data_113;
input 	src_data_114;
input 	src_data_115;
input 	src_data_116;
input 	src_data_86;
input 	Selector5;
input 	Selector12;
input 	src_data_80;
input 	out_data_1;
input 	out_data_0;
input 	Selector6;
input 	Selector13;
input 	src_data_79;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



spw_babasu_altera_merlin_burst_adapter_13_1 \altera_merlin_burst_adapter_13_1.burst_adapter (
	.h2f_ARADDR_0(h2f_ARADDR_0),
	.h2f_ARADDR_1(h2f_ARADDR_1),
	.h2f_ARADDR_2(h2f_ARADDR_2),
	.h2f_ARADDR_3(h2f_ARADDR_3),
	.h2f_ARLEN_0(h2f_ARLEN_0),
	.nxt_in_ready(nxt_in_ready),
	.in_ready_hold1(in_ready_hold),
	.stateST_COMP_TRANS(stateST_COMP_TRANS),
	.out_valid_reg1(out_valid_reg),
	.in_narrow_reg1(in_narrow_reg),
	.in_byteen_reg_3(in_byteen_reg_3),
	.in_byteen_reg_2(in_byteen_reg_2),
	.in_byteen_reg_1(in_byteen_reg_1),
	.in_byteen_reg_0(in_byteen_reg_0),
	.in_data_reg_68(in_data_reg_68),
	.cp_ready(cp_ready),
	.stateST_UNCOMP_WR_SUBBURST(stateST_UNCOMP_WR_SUBBURST),
	.nxt_in_ready1(nxt_in_ready1),
	.sink0_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_116,src_data_115,src_data_114,src_data_113,src_data_112,src_data_111,src_data_110,src_data_109,src_data_108,src_data_107,src_data_106,src_data_105,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_88,src_data_87,
src_data_86,gnd,gnd,gnd,src_data_82,src_data_81,src_data_80,src_data_79,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,saved_grant_1,saved_grant_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_35,src_data_34,src_data_33,
src_data_32,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_payload}),
	.Equal16(Equal16),
	.in_data_reg_0(in_data_reg_0),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_3),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_2),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.Add2(Add2),
	.Add21(Add21),
	.Add22(Add22),
	.Add23(Add23),
	.write_cp_data_77(write_cp_data_77),
	.write_cp_data_78(write_cp_data_78),
	.write_cp_data_75(write_cp_data_75),
	.write_cp_data_74(write_cp_data_74),
	.write_cp_data_76(write_cp_data_76),
	.WideNor0(WideNor0),
	.Equal14(Equal14),
	.nxt_out_eop(nxt_out_eop),
	.src2_valid(src2_valid),
	.src_valid(src_valid),
	.cp_ready1(cp_ready1),
	.in_data_reg_69(in_data_reg_69),
	.src_valid1(src_valid1),
	.out_byte_cnt_reg_2(out_byte_cnt_reg_2),
	.out_uncomp_byte_cnt_reg_5(out_uncomp_byte_cnt_reg_5),
	.out_uncomp_byte_cnt_reg_4(out_uncomp_byte_cnt_reg_4),
	.out_uncomp_byte_cnt_reg_3(out_uncomp_byte_cnt_reg_3),
	.out_uncomp_byte_cnt_reg_2(out_uncomp_byte_cnt_reg_2),
	.out_uncomp_byte_cnt_reg_6(out_uncomp_byte_cnt_reg_6),
	.sink0_endofpacket(src_payload_0),
	.in_data_reg_105(in_data_reg_105),
	.in_data_reg_106(in_data_reg_106),
	.in_data_reg_107(in_data_reg_107),
	.in_data_reg_108(in_data_reg_108),
	.in_data_reg_109(in_data_reg_109),
	.in_data_reg_110(in_data_reg_110),
	.in_data_reg_111(in_data_reg_111),
	.in_data_reg_112(in_data_reg_112),
	.in_data_reg_113(in_data_reg_113),
	.in_data_reg_114(in_data_reg_114),
	.in_data_reg_115(in_data_reg_115),
	.in_data_reg_116(in_data_reg_116),
	.Selector3(Selector3),
	.Selector10(Selector10),
	.base_address_3(base_address_3),
	.Selector4(Selector4),
	.Selector11(Selector11),
	.base_address_2(base_address_2),
	.Selector5(Selector5),
	.Selector12(Selector12),
	.out_data_1(out_data_1),
	.out_data_0(out_data_0),
	.Selector6(Selector6),
	.Selector13(Selector13),
	.clk_clk(clk_clk));

endmodule

module spw_babasu_altera_merlin_burst_adapter_13_1 (
	h2f_ARADDR_0,
	h2f_ARADDR_1,
	h2f_ARADDR_2,
	h2f_ARADDR_3,
	h2f_ARLEN_0,
	nxt_in_ready,
	in_ready_hold1,
	stateST_COMP_TRANS,
	out_valid_reg1,
	in_narrow_reg1,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	in_data_reg_68,
	cp_ready,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready1,
	sink0_data,
	Equal16,
	in_data_reg_0,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	altera_reset_synchronizer_int_chain_out,
	Add2,
	Add21,
	Add22,
	Add23,
	write_cp_data_77,
	write_cp_data_78,
	write_cp_data_75,
	write_cp_data_74,
	write_cp_data_76,
	WideNor0,
	Equal14,
	nxt_out_eop,
	src2_valid,
	src_valid,
	cp_ready1,
	in_data_reg_69,
	src_valid1,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_6,
	sink0_endofpacket,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	Selector3,
	Selector10,
	base_address_3,
	Selector4,
	Selector11,
	base_address_2,
	Selector5,
	Selector12,
	out_data_1,
	out_data_0,
	Selector6,
	Selector13,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARADDR_0;
input 	h2f_ARADDR_1;
input 	h2f_ARADDR_2;
input 	h2f_ARADDR_3;
input 	h2f_ARLEN_0;
output 	nxt_in_ready;
output 	in_ready_hold1;
output 	stateST_COMP_TRANS;
output 	out_valid_reg1;
output 	in_narrow_reg1;
output 	in_byteen_reg_3;
output 	in_byteen_reg_2;
output 	in_byteen_reg_1;
output 	in_byteen_reg_0;
output 	in_data_reg_68;
input 	cp_ready;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready1;
input 	[128:0] sink0_data;
input 	Equal16;
output 	in_data_reg_0;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
input 	altera_reset_synchronizer_int_chain_out;
input 	Add2;
input 	Add21;
input 	Add22;
input 	Add23;
input 	write_cp_data_77;
input 	write_cp_data_78;
input 	write_cp_data_75;
input 	write_cp_data_74;
input 	write_cp_data_76;
input 	WideNor0;
input 	Equal14;
output 	nxt_out_eop;
input 	src2_valid;
input 	src_valid;
input 	cp_ready1;
output 	in_data_reg_69;
input 	src_valid1;
output 	out_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_6;
input 	sink0_endofpacket;
output 	in_data_reg_105;
output 	in_data_reg_106;
output 	in_data_reg_107;
output 	in_data_reg_108;
output 	in_data_reg_109;
output 	in_data_reg_110;
output 	in_data_reg_111;
output 	in_data_reg_112;
output 	in_data_reg_113;
output 	in_data_reg_114;
output 	in_data_reg_115;
output 	in_data_reg_116;
input 	Selector3;
input 	Selector10;
input 	base_address_3;
input 	Selector4;
input 	Selector11;
input 	base_address_2;
input 	Selector5;
input 	Selector12;
input 	out_data_1;
input 	out_data_0;
input 	Selector6;
input 	Selector13;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \align_address_to_size|LessThan0~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt~0_combout ;
wire \Add4~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt[5]~1_combout ;
wire \nxt_uncomp_subburst_byte_cnt[4]~2_combout ;
wire \nxt_uncomp_subburst_byte_cnt[3]~3_combout ;
wire \nxt_uncomp_subburst_byte_cnt[2]~4_combout ;
wire \nxt_uncomp_subburst_byte_cnt[6]~5_combout ;
wire \WideOr0~combout ;
wire \in_valid~combout ;
wire \Selector0~0_combout ;
wire \load_next_out_cmd~combout ;
wire \state.ST_IDLE~q ;
wire \Selector2~0_combout ;
wire \Selector2~1_combout ;
wire \Selector2~2_combout ;
wire \state.ST_UNCOMP_TRANS~q ;
wire \Selector1~0_combout ;
wire \Selector1~1_combout ;
wire \int_bytes_remaining_reg[5]~q ;
wire \d0_int_bytes_remaining[2]~7_combout ;
wire \d0_int_bytes_remaining[2]~8_combout ;
wire \int_bytes_remaining_reg[2]~q ;
wire \d0_int_bytes_remaining[3]~5_combout ;
wire \d0_int_bytes_remaining[3]~6_combout ;
wire \int_bytes_remaining_reg[3]~q ;
wire \Add1~1_combout ;
wire \d0_int_bytes_remaining[4]~4_combout ;
wire \int_bytes_remaining_reg[4]~q ;
wire \Add1~0_combout ;
wire \d0_int_bytes_remaining[5]~0_combout ;
wire \d0_int_bytes_remaining[5]~1_combout ;
wire \int_bytes_remaining_reg[6]~q ;
wire \d0_int_bytes_remaining[6]~2_combout ;
wire \d0_int_bytes_remaining[6]~3_combout ;
wire \new_burst_reg~0_combout ;
wire \new_burst_reg~q ;
wire \WideNor0~0_combout ;
wire \NON_PIPELINED_INPUTS.load_next_cmd~combout ;
wire \in_bytecount_reg_zero~q ;
wire \nxt_out_valid~0_combout ;
wire \LessThan0~0_combout ;
wire \Selector3~0_combout ;
wire \in_size_reg[0]~q ;
wire \in_size_reg[2]~q ;
wire \in_size_reg[1]~q ;
wire \ShiftLeft0~0_combout ;
wire \ShiftLeft0~1_combout ;
wire \int_byte_cnt_narrow_reg[3]~q ;
wire \ShiftLeft0~2_combout ;
wire \int_byte_cnt_narrow_reg[2]~q ;
wire \ShiftLeft0~3_combout ;
wire \ShiftLeft0~4_combout ;
wire \int_byte_cnt_narrow_reg[1]~q ;
wire \int_byte_cnt_narrow_reg[0]~q ;
wire \Add0~13_sumout ;
wire \d0_int_nxt_addr[0]~3_combout ;
wire \in_burstwrap_reg[0]~q ;
wire \nxt_addr[0]~0_combout ;
wire \int_nxt_addr_reg[0]~q ;
wire \d0_int_nxt_addr[0]~4_combout ;
wire \int_nxt_addr_reg_dly[0]~q ;
wire \Add0~14 ;
wire \Add0~9_sumout ;
wire \in_burstwrap_reg[1]~q ;
wire \nxt_addr[1]~4_combout ;
wire \int_nxt_addr_reg[1]~q ;
wire \d0_int_nxt_addr[1]~7_combout ;
wire \d0_int_nxt_addr[1]~2_combout ;
wire \int_nxt_addr_reg_dly[1]~q ;
wire \Add0~10 ;
wire \Add0~6 ;
wire \Add0~1_sumout ;
wire \in_burstwrap_reg[3]~q ;
wire \nxt_addr[3]~12_combout ;
wire \int_nxt_addr_reg[3]~q ;
wire \d0_int_nxt_addr[3]~5_combout ;
wire \d0_int_nxt_addr[3]~0_combout ;
wire \Add0~5_sumout ;
wire \in_burstwrap_reg[2]~q ;
wire \nxt_addr[2]~8_combout ;
wire \int_nxt_addr_reg[2]~q ;
wire \d0_int_nxt_addr[2]~6_combout ;
wire \d0_int_nxt_addr[2]~1_combout ;
wire \in_eop_reg~q ;


spw_babasu_altera_merlin_address_alignment_1 align_address_to_size(
	.new_burst_reg(\new_burst_reg~q ),
	.src_data_86(sink0_data[86]),
	.in_size_reg_0(\in_size_reg[0]~q ),
	.ShiftLeft0(\ShiftLeft0~3_combout ),
	.LessThan0(\align_address_to_size|LessThan0~0_combout ));

cyclonev_lcell_comb \nxt_in_ready~1 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!in_ready_hold1),
	.datac(!out_valid_reg1),
	.datad(!cp_ready),
	.datae(!stateST_COMP_TRANS),
	.dataf(!\new_burst_reg~q ),
	.datag(!stateST_UNCOMP_WR_SUBBURST),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~1 .extended_lut = "on";
defparam \nxt_in_ready~1 .lut_mask = 64'h2020F0F02020F0FF;
defparam \nxt_in_ready~1 .shared_arith = "off";

dffeas in_ready_hold(
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(in_ready_hold1),
	.prn(vcc));
defparam in_ready_hold.is_wysiwyg = "true";
defparam in_ready_hold.power_up = "low";

dffeas \state.ST_COMP_TRANS (
	.clk(clk_clk),
	.d(\Selector1~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_COMP_TRANS),
	.prn(vcc));
defparam \state.ST_COMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_COMP_TRANS .power_up = "low";

dffeas out_valid_reg(
	.clk(clk_clk),
	.d(\nxt_out_valid~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_valid_reg1),
	.prn(vcc));
defparam out_valid_reg.is_wysiwyg = "true";
defparam out_valid_reg.power_up = "low";

dffeas in_narrow_reg(
	.clk(clk_clk),
	.d(\LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_narrow_reg1),
	.prn(vcc));
defparam in_narrow_reg.is_wysiwyg = "true";
defparam in_narrow_reg.power_up = "low";

dffeas \in_byteen_reg[3] (
	.clk(clk_clk),
	.d(sink0_data[35]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_3),
	.prn(vcc));
defparam \in_byteen_reg[3] .is_wysiwyg = "true";
defparam \in_byteen_reg[3] .power_up = "low";

dffeas \in_byteen_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[34]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_2),
	.prn(vcc));
defparam \in_byteen_reg[2] .is_wysiwyg = "true";
defparam \in_byteen_reg[2] .power_up = "low";

dffeas \in_byteen_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[33]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_1),
	.prn(vcc));
defparam \in_byteen_reg[1] .is_wysiwyg = "true";
defparam \in_byteen_reg[1] .power_up = "low";

dffeas \in_byteen_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[32]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_0),
	.prn(vcc));
defparam \in_byteen_reg[0] .is_wysiwyg = "true";
defparam \in_byteen_reg[0] .power_up = "low";

dffeas \in_data_reg[68] (
	.clk(clk_clk),
	.d(sink0_data[68]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_68),
	.prn(vcc));
defparam \in_data_reg[68] .is_wysiwyg = "true";
defparam \in_data_reg[68] .power_up = "low";

dffeas \state.ST_UNCOMP_WR_SUBBURST (
	.clk(clk_clk),
	.d(\Selector3~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_UNCOMP_WR_SUBBURST),
	.prn(vcc));
defparam \state.ST_UNCOMP_WR_SUBBURST .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_WR_SUBBURST .power_up = "low";

cyclonev_lcell_comb \nxt_in_ready~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!out_valid_reg1),
	.datac(!cp_ready),
	.datad(!\state.ST_UNCOMP_TRANS~q ),
	.datae(!stateST_UNCOMP_WR_SUBBURST),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~0 .extended_lut = "off";
defparam \nxt_in_ready~0 .lut_mask = 64'h008A8A8A008A8A8A;
defparam \nxt_in_ready~0 .shared_arith = "off";

dffeas \in_data_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[0]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_0),
	.prn(vcc));
defparam \in_data_reg[0] .is_wysiwyg = "true";
defparam \in_data_reg[0] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[3] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[3]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_3),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[3] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[2] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[2]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_2),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[2] .power_up = "low";

cyclonev_lcell_comb \nxt_out_eop~0 (
	.dataa(!\in_eop_reg~q ),
	.datab(!stateST_COMP_TRANS),
	.datac(!\new_burst_reg~q ),
	.datad(!cp_ready),
	.datae(!\in_bytecount_reg_zero~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_out_eop),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_eop~0 .extended_lut = "off";
defparam \nxt_out_eop~0 .lut_mask = 64'h4447774744477747;
defparam \nxt_out_eop~0 .shared_arith = "off";

dffeas \in_data_reg[69] (
	.clk(clk_clk),
	.d(sink0_data[69]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_69),
	.prn(vcc));
defparam \in_data_reg[69] .is_wysiwyg = "true";
defparam \in_data_reg[69] .power_up = "low";

dffeas \out_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[5] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[5]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_5),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[5] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[5] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[4] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[4]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_4),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[4] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[4] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[3] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[3]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_3),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[3] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[3] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[2]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[6] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[6]~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_6),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[6] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[6] .power_up = "low";

dffeas \in_data_reg[105] (
	.clk(clk_clk),
	.d(sink0_data[105]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_105),
	.prn(vcc));
defparam \in_data_reg[105] .is_wysiwyg = "true";
defparam \in_data_reg[105] .power_up = "low";

dffeas \in_data_reg[106] (
	.clk(clk_clk),
	.d(sink0_data[106]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_106),
	.prn(vcc));
defparam \in_data_reg[106] .is_wysiwyg = "true";
defparam \in_data_reg[106] .power_up = "low";

dffeas \in_data_reg[107] (
	.clk(clk_clk),
	.d(sink0_data[107]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_107),
	.prn(vcc));
defparam \in_data_reg[107] .is_wysiwyg = "true";
defparam \in_data_reg[107] .power_up = "low";

dffeas \in_data_reg[108] (
	.clk(clk_clk),
	.d(sink0_data[108]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_108),
	.prn(vcc));
defparam \in_data_reg[108] .is_wysiwyg = "true";
defparam \in_data_reg[108] .power_up = "low";

dffeas \in_data_reg[109] (
	.clk(clk_clk),
	.d(sink0_data[109]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_109),
	.prn(vcc));
defparam \in_data_reg[109] .is_wysiwyg = "true";
defparam \in_data_reg[109] .power_up = "low";

dffeas \in_data_reg[110] (
	.clk(clk_clk),
	.d(sink0_data[110]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_110),
	.prn(vcc));
defparam \in_data_reg[110] .is_wysiwyg = "true";
defparam \in_data_reg[110] .power_up = "low";

dffeas \in_data_reg[111] (
	.clk(clk_clk),
	.d(sink0_data[111]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_111),
	.prn(vcc));
defparam \in_data_reg[111] .is_wysiwyg = "true";
defparam \in_data_reg[111] .power_up = "low";

dffeas \in_data_reg[112] (
	.clk(clk_clk),
	.d(sink0_data[112]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_112),
	.prn(vcc));
defparam \in_data_reg[112] .is_wysiwyg = "true";
defparam \in_data_reg[112] .power_up = "low";

dffeas \in_data_reg[113] (
	.clk(clk_clk),
	.d(sink0_data[113]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_113),
	.prn(vcc));
defparam \in_data_reg[113] .is_wysiwyg = "true";
defparam \in_data_reg[113] .power_up = "low";

dffeas \in_data_reg[114] (
	.clk(clk_clk),
	.d(sink0_data[114]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_114),
	.prn(vcc));
defparam \in_data_reg[114] .is_wysiwyg = "true";
defparam \in_data_reg[114] .power_up = "low";

dffeas \in_data_reg[115] (
	.clk(clk_clk),
	.d(sink0_data[115]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_115),
	.prn(vcc));
defparam \in_data_reg[115] .is_wysiwyg = "true";
defparam \in_data_reg[115] .power_up = "low";

dffeas \in_data_reg[116] (
	.clk(clk_clk),
	.d(sink0_data[116]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_116),
	.prn(vcc));
defparam \in_data_reg[116] .is_wysiwyg = "true";
defparam \in_data_reg[116] .power_up = "low";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt~0 (
	.dataa(!out_valid_reg1),
	.datab(!cp_ready),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt~0 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt~0 .lut_mask = 64'h1111111111111111;
defparam \nxt_uncomp_subburst_byte_cnt~0 .shared_arith = "off";

cyclonev_lcell_comb \Add4~0 (
	.dataa(!out_uncomp_byte_cnt_reg_4),
	.datab(!out_uncomp_byte_cnt_reg_3),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add4~0 .extended_lut = "off";
defparam \Add4~0 .lut_mask = 64'h0800080008000800;
defparam \Add4~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[5]~1 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!\Add4~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[5]~1 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[5]~1 .lut_mask = 64'h0F4EA5E40F4EA5E4;
defparam \nxt_uncomp_subburst_byte_cnt[5]~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[4]~2 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!out_uncomp_byte_cnt_reg_3),
	.datae(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.dataf(!out_uncomp_byte_cnt_reg_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[4]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[4]~2 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[4]~2 .lut_mask = 64'h0F0FE44E0F0F4E4E;
defparam \nxt_uncomp_subburst_byte_cnt[4]~2 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[3]~3 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!out_uncomp_byte_cnt_reg_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[3]~3 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[3]~3 .lut_mask = 64'h0FE40F4E0FE40F4E;
defparam \nxt_uncomp_subburst_byte_cnt[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[2]~4 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[2]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[2]~4 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[2]~4 .lut_mask = 64'h0EF40EF40EF40EF4;
defparam \nxt_uncomp_subburst_byte_cnt[2]~4 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[6]~5 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!\Add4~0_combout ),
	.dataf(!out_uncomp_byte_cnt_reg_6),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[6]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[6]~5 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[6]~5 .lut_mask = 64'h0044A0E4FFEE5F4E;
defparam \nxt_uncomp_subburst_byte_cnt[6]~5 .shared_arith = "off";

cyclonev_lcell_comb WideOr0(
	.dataa(!\nxt_uncomp_subburst_byte_cnt[5]~1_combout ),
	.datab(!\nxt_uncomp_subburst_byte_cnt[4]~2_combout ),
	.datac(!\nxt_uncomp_subburst_byte_cnt[3]~3_combout ),
	.datad(!\nxt_uncomp_subburst_byte_cnt[2]~4_combout ),
	.datae(!\nxt_uncomp_subburst_byte_cnt[6]~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr0.extended_lut = "off";
defparam WideOr0.lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam WideOr0.shared_arith = "off";

cyclonev_lcell_comb in_valid(
	.dataa(!in_ready_hold1),
	.datab(!Equal16),
	.datac(!Equal14),
	.datad(!sink0_data[68]),
	.datae(!src2_valid),
	.dataf(!src_valid),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\in_valid~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam in_valid.extended_lut = "off";
defparam in_valid.lut_mask = 64'h0000000155555555;
defparam in_valid.shared_arith = "off";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!sink0_data[69]),
	.datab(!nxt_out_eop),
	.datac(!sink0_data[68]),
	.datad(!\in_valid~combout ),
	.datae(!\state.ST_IDLE~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'h005FCCFF005FCCFF;
defparam \Selector0~0 .shared_arith = "off";

cyclonev_lcell_comb load_next_out_cmd(
	.dataa(!out_valid_reg1),
	.datab(!cp_ready),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\load_next_out_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam load_next_out_cmd.extended_lut = "off";
defparam load_next_out_cmd.lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam load_next_out_cmd.shared_arith = "off";

dffeas \state.ST_IDLE (
	.clk(clk_clk),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_IDLE~q ),
	.prn(vcc));
defparam \state.ST_IDLE .is_wysiwyg = "true";
defparam \state.ST_IDLE .power_up = "low";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!nxt_out_eop),
	.datac(!stateST_UNCOMP_WR_SUBBURST),
	.datad(!\state.ST_IDLE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'h00EC00EC00EC00EC;
defparam \Selector2~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~1 (
	.dataa(!in_ready_hold1),
	.datab(!Equal16),
	.datac(!Equal14),
	.datad(!sink0_data[68]),
	.datae(!src2_valid),
	.dataf(!\Selector2~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~1 .extended_lut = "off";
defparam \Selector2~1 .lut_mask = 64'h0000000100000000;
defparam \Selector2~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~2 (
	.dataa(!\WideOr0~combout ),
	.datab(!\Selector2~1_combout ),
	.datac(!\in_valid~combout ),
	.datad(!nxt_out_eop),
	.datae(!\state.ST_UNCOMP_TRANS~q ),
	.dataf(!sink0_data[69]),
	.datag(!stateST_UNCOMP_WR_SUBBURST),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~2 .extended_lut = "on";
defparam \Selector2~2 .lut_mask = 64'h3B33BB3F0A00AA00;
defparam \Selector2~2 .shared_arith = "off";

dffeas \state.ST_UNCOMP_TRANS (
	.clk(clk_clk),
	.d(\Selector2~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_UNCOMP_TRANS~q ),
	.prn(vcc));
defparam \state.ST_UNCOMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_TRANS .power_up = "low";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!nxt_out_eop),
	.datac(!\state.ST_UNCOMP_TRANS~q ),
	.datad(!stateST_UNCOMP_WR_SUBBURST),
	.datae(!\state.ST_IDLE~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'h0000A8880000A888;
defparam \Selector1~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~1 (
	.dataa(!sink0_data[69]),
	.datab(!stateST_COMP_TRANS),
	.datac(!nxt_out_eop),
	.datad(!sink0_data[68]),
	.datae(!\in_valid~combout ),
	.dataf(!\Selector1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~1 .extended_lut = "off";
defparam \Selector1~1 .lut_mask = 64'h3030777530303330;
defparam \Selector1~1 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[5] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[5]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[5]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[5] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[5] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[2]~7 (
	.dataa(!h2f_ARLEN_0),
	.datab(!sink0_data[69]),
	.datac(!sink0_data[68]),
	.datad(!write_cp_data_74),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[2]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[2]~7 .extended_lut = "off";
defparam \d0_int_bytes_remaining[2]~7 .lut_mask = 64'h2F222F222F222F22;
defparam \d0_int_bytes_remaining[2]~7 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[2]~8 (
	.dataa(!\new_burst_reg~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\int_bytes_remaining_reg[2]~q ),
	.datad(!\d0_int_bytes_remaining[2]~7_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[2]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[2]~8 .extended_lut = "off";
defparam \d0_int_bytes_remaining[2]~8 .lut_mask = 64'h287D287D287D287D;
defparam \d0_int_bytes_remaining[2]~8 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[2] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[2]~8_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[2]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[2] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[3]~5 (
	.dataa(!sink0_data[69]),
	.datab(!sink0_data[68]),
	.datac(!write_cp_data_75),
	.datad(!Add2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[3]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[3]~5 .extended_lut = "off";
defparam \d0_int_bytes_remaining[3]~5 .lut_mask = 64'h0357035703570357;
defparam \d0_int_bytes_remaining[3]~5 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[3]~6 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\int_bytes_remaining_reg[3]~q ),
	.datac(!out_byte_cnt_reg_2),
	.datad(!\int_bytes_remaining_reg[2]~q ),
	.datae(!\d0_int_bytes_remaining[3]~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[3]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[3]~6 .extended_lut = "off";
defparam \d0_int_bytes_remaining[3]~6 .lut_mask = 64'h28227D7728227D77;
defparam \d0_int_bytes_remaining[3]~6 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[3] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[3]~6_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[3]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[3] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[3] .power_up = "low";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!\int_bytes_remaining_reg[4]~q ),
	.datab(!\int_bytes_remaining_reg[3]~q ),
	.datac(!out_byte_cnt_reg_2),
	.datad(!\int_bytes_remaining_reg[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'hA6AAA6AAA6AAA6AA;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[4]~4 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!sink0_data[68]),
	.datad(!write_cp_data_76),
	.datae(!Add21),
	.dataf(!\Add1~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[4]~4 .extended_lut = "off";
defparam \d0_int_bytes_remaining[4]~4 .lut_mask = 64'hCCCFDDDF00031113;
defparam \d0_int_bytes_remaining[4]~4 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[4] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[4]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[4]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[4] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[4] .power_up = "low";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!\int_bytes_remaining_reg[4]~q ),
	.datab(!\int_bytes_remaining_reg[3]~q ),
	.datac(!out_byte_cnt_reg_2),
	.datad(!\int_bytes_remaining_reg[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h0800080008000800;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[5]~0 (
	.dataa(!sink0_data[69]),
	.datab(!sink0_data[68]),
	.datac(!write_cp_data_77),
	.datad(!Add22),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[5]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[5]~0 .extended_lut = "off";
defparam \d0_int_bytes_remaining[5]~0 .lut_mask = 64'h0357035703570357;
defparam \d0_int_bytes_remaining[5]~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[5]~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\int_bytes_remaining_reg[5]~q ),
	.datac(!\Add1~0_combout ),
	.datad(!\d0_int_bytes_remaining[5]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[5]~1 .extended_lut = "off";
defparam \d0_int_bytes_remaining[5]~1 .lut_mask = 64'h287D287D287D287D;
defparam \d0_int_bytes_remaining[5]~1 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[6] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[6]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[6]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[6] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[6] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[6]~2 (
	.dataa(!sink0_data[69]),
	.datab(!sink0_data[68]),
	.datac(!write_cp_data_78),
	.datad(!Add23),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[6]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[6]~2 .extended_lut = "off";
defparam \d0_int_bytes_remaining[6]~2 .lut_mask = 64'h0357035703570357;
defparam \d0_int_bytes_remaining[6]~2 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[6]~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\int_bytes_remaining_reg[5]~q ),
	.datac(!\Add1~0_combout ),
	.datad(!\int_bytes_remaining_reg[6]~q ),
	.datae(!\d0_int_bytes_remaining[6]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[6]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[6]~3 .extended_lut = "off";
defparam \d0_int_bytes_remaining[6]~3 .lut_mask = 64'h08A25DF708A25DF7;
defparam \d0_int_bytes_remaining[6]~3 .shared_arith = "off";

cyclonev_lcell_comb \new_burst_reg~0 (
	.dataa(!\Selector1~1_combout ),
	.datab(!\d0_int_bytes_remaining[5]~1_combout ),
	.datac(!\d0_int_bytes_remaining[6]~3_combout ),
	.datad(!\d0_int_bytes_remaining[4]~4_combout ),
	.datae(!\d0_int_bytes_remaining[3]~6_combout ),
	.dataf(!\d0_int_bytes_remaining[2]~8_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\new_burst_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \new_burst_reg~0 .extended_lut = "off";
defparam \new_burst_reg~0 .lut_mask = 64'hAAAAAAAAEAAAAAAA;
defparam \new_burst_reg~0 .shared_arith = "off";

dffeas new_burst_reg(
	.clk(clk_clk),
	.d(\new_burst_reg~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\new_burst_reg~q ),
	.prn(vcc));
defparam new_burst_reg.is_wysiwyg = "true";
defparam new_burst_reg.power_up = "low";

cyclonev_lcell_comb \WideNor0~0 (
	.dataa(!sink0_data[69]),
	.datab(!sink0_data[68]),
	.datac(!WideNor0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideNor0~0 .extended_lut = "off";
defparam \WideNor0~0 .lut_mask = 64'h8A8A8A8A8A8A8A8A;
defparam \WideNor0~0 .shared_arith = "off";

cyclonev_lcell_comb \NON_PIPELINED_INPUTS.load_next_cmd (
	.dataa(!in_ready_hold1),
	.datab(!nxt_in_ready1),
	.datac(!nxt_in_ready),
	.datad(!src_valid),
	.datae(!src_valid1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \NON_PIPELINED_INPUTS.load_next_cmd .extended_lut = "off";
defparam \NON_PIPELINED_INPUTS.load_next_cmd .lut_mask = 64'h0015151500151515;
defparam \NON_PIPELINED_INPUTS.load_next_cmd .shared_arith = "off";

dffeas in_bytecount_reg_zero(
	.clk(clk_clk),
	.d(\WideNor0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_bytecount_reg_zero~q ),
	.prn(vcc));
defparam in_bytecount_reg_zero.is_wysiwyg = "true";
defparam in_bytecount_reg_zero.power_up = "low";

cyclonev_lcell_comb \nxt_out_valid~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!\new_burst_reg~q ),
	.datac(!\in_bytecount_reg_zero~q ),
	.datad(!\in_valid~combout ),
	.datae(!cp_ready1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_valid~0 .extended_lut = "off";
defparam \nxt_out_valid~0 .lut_mask = 64'h50FF44FF50FF44FF;
defparam \nxt_out_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!sink0_data[87]),
	.datab(!sink0_data[88]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h8888888888888888;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~0 (
	.dataa(!nxt_out_eop),
	.datab(!\state.ST_UNCOMP_TRANS~q ),
	.datac(!stateST_UNCOMP_WR_SUBBURST),
	.datad(!\WideOr0~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'h002A002A002A002A;
defparam \Selector3~0 .shared_arith = "off";

dffeas \in_size_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[86]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[0]~q ),
	.prn(vcc));
defparam \in_size_reg[0] .is_wysiwyg = "true";
defparam \in_size_reg[0] .power_up = "low";

dffeas \in_size_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[88]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[2]~q ),
	.prn(vcc));
defparam \in_size_reg[2] .is_wysiwyg = "true";
defparam \in_size_reg[2] .power_up = "low";

dffeas \in_size_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[87]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[1]~q ),
	.prn(vcc));
defparam \in_size_reg[1] .is_wysiwyg = "true";
defparam \in_size_reg[1] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[87]),
	.datac(!sink0_data[88]),
	.datad(!\in_size_reg[2]~q ),
	.datae(!\in_size_reg[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~0 .extended_lut = "off";
defparam \ShiftLeft0~0 .lut_mask = 64'h1010BA101010BA10;
defparam \ShiftLeft0~0 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~1 .extended_lut = "off";
defparam \ShiftLeft0~1 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~1 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[3] (
	.clk(clk_clk),
	.d(\ShiftLeft0~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[3]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[3] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[3] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~2 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~2 .extended_lut = "off";
defparam \ShiftLeft0~2 .lut_mask = 64'h00E400E400E400E4;
defparam \ShiftLeft0~2 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[2] (
	.clk(clk_clk),
	.d(\ShiftLeft0~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[2]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[2] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[2] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[87]),
	.datac(!sink0_data[88]),
	.datad(!\in_size_reg[2]~q ),
	.datae(!\in_size_reg[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~3 .extended_lut = "off";
defparam \ShiftLeft0~3 .lut_mask = 64'hEA404040EA404040;
defparam \ShiftLeft0~3 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~4 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~4 .extended_lut = "off";
defparam \ShiftLeft0~4 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~4 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[1] (
	.clk(clk_clk),
	.d(\ShiftLeft0~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[1]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[1] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[1] .power_up = "low";

dffeas \int_byte_cnt_narrow_reg[0] (
	.clk(clk_clk),
	.d(\align_address_to_size|LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[0]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[0] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[0] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[0]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~3 (
	.dataa(!h2f_ARADDR_0),
	.datab(!sink0_data[69]),
	.datac(!sink0_data[68]),
	.datad(!out_data_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~3 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~3 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[0]~3 .shared_arith = "off";

dffeas \in_burstwrap_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[79]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[0]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[0] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[0] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[0]~0 (
	.dataa(!Selector13),
	.datab(!Selector6),
	.datac(!sink0_data[68]),
	.datad(!sink0_data[69]),
	.datae(!\new_burst_reg~q ),
	.dataf(!\d0_int_nxt_addr[0]~4_combout ),
	.datag(!\in_burstwrap_reg[0]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[0]~0 .extended_lut = "on";
defparam \nxt_addr[0]~0 .lut_mask = 64'h00000000F0F0FCA8;
defparam \nxt_addr[0]~0 .shared_arith = "off";

dffeas \int_nxt_addr_reg[0] (
	.clk(clk_clk),
	.d(\nxt_addr[0]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[0] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~4 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\Add0~13_sumout ),
	.datac(!\align_address_to_size|LessThan0~0_combout ),
	.datad(!\d0_int_nxt_addr[0]~3_combout ),
	.datae(!\int_nxt_addr_reg[0]~q ),
	.dataf(!\in_burstwrap_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~4 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~4 .lut_mask = 64'h0005AAAF2227AAAF;
defparam \d0_int_nxt_addr[0]~4 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[0] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[0]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[0] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[1]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[1]~q ),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \in_burstwrap_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[80]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[1]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[1] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[1] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[1]~4 (
	.dataa(!Selector12),
	.datab(!Selector5),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!\new_burst_reg~q ),
	.dataf(!\d0_int_nxt_addr[1]~2_combout ),
	.datag(!\in_burstwrap_reg[1]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[1]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[1]~4 .extended_lut = "on";
defparam \nxt_addr[1]~4 .lut_mask = 64'h00000000F0F0FAC8;
defparam \nxt_addr[1]~4 .shared_arith = "off";

dffeas \int_nxt_addr_reg[1] (
	.clk(clk_clk),
	.d(\nxt_addr[1]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[1] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~7 (
	.dataa(!h2f_ARADDR_1),
	.datab(!sink0_data[69]),
	.datac(!sink0_data[68]),
	.datad(!out_data_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~7 .extended_lut = "off";
defparam \d0_int_nxt_addr[1]~7 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[1]~7 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~2 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\Add0~9_sumout ),
	.datac(!\in_burstwrap_reg[1]~q ),
	.datad(!\int_nxt_addr_reg[1]~q ),
	.datae(!\ShiftLeft0~3_combout ),
	.dataf(!\d0_int_nxt_addr[1]~7_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~2 .extended_lut = "off";
defparam \d0_int_nxt_addr[1]~2 .lut_mask = 64'h02AA02AA02AA57FF;
defparam \d0_int_nxt_addr[1]~2 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[1] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[1]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[1] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_2),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[2]~q ),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[3]~q ),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

dffeas \in_burstwrap_reg[3] (
	.clk(clk_clk),
	.d(sink0_data[82]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[3]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[3] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[3] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[3]~12 (
	.dataa(!Selector10),
	.datab(!Selector3),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!\new_burst_reg~q ),
	.dataf(!\d0_int_nxt_addr[3]~0_combout ),
	.datag(!\in_burstwrap_reg[3]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[3]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[3]~12 .extended_lut = "on";
defparam \nxt_addr[3]~12 .lut_mask = 64'h00000000F0F0FAC8;
defparam \nxt_addr[3]~12 .shared_arith = "off";

dffeas \int_nxt_addr_reg[3] (
	.clk(clk_clk),
	.d(\nxt_addr[3]~12_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[3]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[3] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~5 (
	.dataa(!\Add0~1_sumout ),
	.datab(!\in_burstwrap_reg[3]~q ),
	.datac(!\int_nxt_addr_reg[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~5 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~5 .lut_mask = 64'hE0E0E0E0E0E0E0E0;
defparam \d0_int_nxt_addr[3]~5 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!h2f_ARADDR_3),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!base_address_3),
	.dataf(!\d0_int_nxt_addr[3]~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~0 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~0 .lut_mask = 64'hABABABFF01010155;
defparam \d0_int_nxt_addr[3]~0 .shared_arith = "off";

dffeas \in_burstwrap_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[81]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[2]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[2] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[2] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[2]~8 (
	.dataa(!Selector11),
	.datab(!Selector4),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!\new_burst_reg~q ),
	.dataf(!\d0_int_nxt_addr[2]~1_combout ),
	.datag(!\in_burstwrap_reg[2]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[2]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[2]~8 .extended_lut = "on";
defparam \nxt_addr[2]~8 .lut_mask = 64'h00000000F0F0FAC8;
defparam \nxt_addr[2]~8 .shared_arith = "off";

dffeas \int_nxt_addr_reg[2] (
	.clk(clk_clk),
	.d(\nxt_addr[2]~8_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[2]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~6 (
	.dataa(!\Add0~5_sumout ),
	.datab(!\in_burstwrap_reg[2]~q ),
	.datac(!\int_nxt_addr_reg[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~6 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~6 .lut_mask = 64'hE0E0E0E0E0E0E0E0;
defparam \d0_int_nxt_addr[2]~6 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!h2f_ARADDR_2),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!base_address_2),
	.dataf(!\d0_int_nxt_addr[2]~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~1 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~1 .lut_mask = 64'hABABABFF01010155;
defparam \d0_int_nxt_addr[2]~1 .shared_arith = "off";

dffeas in_eop_reg(
	.clk(clk_clk),
	.d(sink0_endofpacket),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_eop_reg~q ),
	.prn(vcc));
defparam in_eop_reg.is_wysiwyg = "true";
defparam in_eop_reg.power_up = "low";

endmodule

module spw_babasu_altera_merlin_address_alignment_1 (
	new_burst_reg,
	src_data_86,
	in_size_reg_0,
	ShiftLeft0,
	LessThan0)/* synthesis synthesis_greybox=0 */;
input 	new_burst_reg;
input 	src_data_86;
input 	in_size_reg_0;
input 	ShiftLeft0;
output 	LessThan0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!new_burst_reg),
	.datab(!src_data_86),
	.datac(!in_size_reg_0),
	.datad(!ShiftLeft0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan0),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h00E400E400E400E4;
defparam \LessThan0~0 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_burst_adapter_1 (
	h2f_ARADDR_0,
	h2f_ARADDR_1,
	h2f_ARADDR_2,
	h2f_ARADDR_3,
	h2f_ARBURST_0,
	h2f_ARBURST_1,
	h2f_ARID_0,
	h2f_ARID_1,
	h2f_ARID_2,
	h2f_ARID_3,
	h2f_ARID_4,
	h2f_ARID_5,
	h2f_ARID_6,
	h2f_ARID_7,
	h2f_ARID_8,
	h2f_ARID_9,
	h2f_ARID_10,
	h2f_ARID_11,
	h2f_ARLEN_0,
	Add5,
	Add51,
	in_ready_hold,
	saved_grant_1,
	stateST_COMP_TRANS,
	mem_used_1,
	in_data_reg_69,
	in_narrow_reg,
	cp_ready,
	cp_ready1,
	nxt_out_eop,
	out_valid_reg,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready,
	altera_reset_synchronizer_int_chain_out,
	Decoder1,
	Add2,
	Add21,
	Add22,
	Add23,
	nxt_in_ready1,
	src_valid,
	out_byte_cnt_reg_2,
	cp_ready2,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_6,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	Selector10,
	Selector101,
	Selector11,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	Selector12,
	src_payload,
	src_payload1,
	src_payload2,
	Selector13,
	nxt_out_burstwrap_1,
	nxt_addr_2,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARADDR_0;
input 	h2f_ARADDR_1;
input 	h2f_ARADDR_2;
input 	h2f_ARADDR_3;
input 	h2f_ARBURST_0;
input 	h2f_ARBURST_1;
input 	h2f_ARID_0;
input 	h2f_ARID_1;
input 	h2f_ARID_2;
input 	h2f_ARID_3;
input 	h2f_ARID_4;
input 	h2f_ARID_5;
input 	h2f_ARID_6;
input 	h2f_ARID_7;
input 	h2f_ARID_8;
input 	h2f_ARID_9;
input 	h2f_ARID_10;
input 	h2f_ARID_11;
input 	h2f_ARLEN_0;
input 	Add5;
input 	Add51;
input 	in_ready_hold;
input 	saved_grant_1;
output 	stateST_COMP_TRANS;
input 	mem_used_1;
output 	in_data_reg_69;
output 	in_narrow_reg;
input 	cp_ready;
input 	cp_ready1;
output 	nxt_out_eop;
output 	out_valid_reg;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready;
input 	altera_reset_synchronizer_int_chain_out;
input 	Decoder1;
input 	Add2;
input 	Add21;
input 	Add22;
input 	Add23;
output 	nxt_in_ready1;
input 	src_valid;
output 	out_byte_cnt_reg_2;
input 	cp_ready2;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_6;
output 	in_data_reg_105;
output 	in_data_reg_106;
output 	in_data_reg_107;
output 	in_data_reg_108;
output 	in_data_reg_109;
output 	in_data_reg_110;
output 	in_data_reg_111;
output 	in_data_reg_112;
output 	in_data_reg_113;
output 	in_data_reg_114;
output 	in_data_reg_115;
output 	in_data_reg_116;
input 	Selector10;
input 	Selector101;
input 	Selector11;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
input 	Selector12;
input 	src_payload;
input 	src_payload1;
input 	src_payload2;
input 	Selector13;
input 	nxt_out_burstwrap_1;
input 	nxt_addr_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



spw_babasu_altera_merlin_burst_adapter_13_1_1 \altera_merlin_burst_adapter_13_1.burst_adapter (
	.h2f_ARADDR_0(h2f_ARADDR_0),
	.h2f_ARADDR_1(h2f_ARADDR_1),
	.h2f_ARADDR_2(h2f_ARADDR_2),
	.h2f_ARADDR_3(h2f_ARADDR_3),
	.h2f_ARBURST_0(h2f_ARBURST_0),
	.h2f_ARBURST_1(h2f_ARBURST_1),
	.sink0_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,h2f_ARID_11,h2f_ARID_10,h2f_ARID_9,h2f_ARID_8,h2f_ARID_7,h2f_ARID_6,h2f_ARID_5,h2f_ARID_4,h2f_ARID_3,h2f_ARID_2,h2f_ARID_1,h2f_ARID_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_payload1,src_payload2,src_payload,gnd,gnd,gnd,
Selector101,Selector11,Selector12,Selector13,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,saved_grant_1,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.h2f_ARLEN_0(h2f_ARLEN_0),
	.Add5(Add5),
	.Add51(Add51),
	.in_ready_hold(in_ready_hold),
	.stateST_COMP_TRANS(stateST_COMP_TRANS),
	.mem_used_1(mem_used_1),
	.in_data_reg_69(in_data_reg_69),
	.in_narrow_reg1(in_narrow_reg),
	.cp_ready(cp_ready),
	.cp_ready1(cp_ready1),
	.nxt_out_eop(nxt_out_eop),
	.out_valid_reg1(out_valid_reg),
	.stateST_UNCOMP_WR_SUBBURST(stateST_UNCOMP_WR_SUBBURST),
	.nxt_in_ready(nxt_in_ready),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.Decoder1(Decoder1),
	.Add2(Add2),
	.Add21(Add21),
	.Add22(Add22),
	.Add23(Add23),
	.nxt_in_ready1(nxt_in_ready1),
	.src_valid(src_valid),
	.out_byte_cnt_reg_2(out_byte_cnt_reg_2),
	.cp_ready2(cp_ready2),
	.out_uncomp_byte_cnt_reg_3(out_uncomp_byte_cnt_reg_3),
	.out_uncomp_byte_cnt_reg_2(out_uncomp_byte_cnt_reg_2),
	.out_uncomp_byte_cnt_reg_4(out_uncomp_byte_cnt_reg_4),
	.out_uncomp_byte_cnt_reg_5(out_uncomp_byte_cnt_reg_5),
	.out_uncomp_byte_cnt_reg_6(out_uncomp_byte_cnt_reg_6),
	.in_data_reg_105(in_data_reg_105),
	.in_data_reg_106(in_data_reg_106),
	.in_data_reg_107(in_data_reg_107),
	.in_data_reg_108(in_data_reg_108),
	.in_data_reg_109(in_data_reg_109),
	.in_data_reg_110(in_data_reg_110),
	.in_data_reg_111(in_data_reg_111),
	.in_data_reg_112(in_data_reg_112),
	.in_data_reg_113(in_data_reg_113),
	.in_data_reg_114(in_data_reg_114),
	.in_data_reg_115(in_data_reg_115),
	.in_data_reg_116(in_data_reg_116),
	.Selector10(Selector10),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_3),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_2),
	.nxt_out_burstwrap_1(nxt_out_burstwrap_1),
	.nxt_addr_2(nxt_addr_2),
	.clk_clk(clk_clk));

endmodule

module spw_babasu_altera_merlin_burst_adapter_13_1_1 (
	h2f_ARADDR_0,
	h2f_ARADDR_1,
	h2f_ARADDR_2,
	h2f_ARADDR_3,
	h2f_ARBURST_0,
	h2f_ARBURST_1,
	sink0_data,
	h2f_ARLEN_0,
	Add5,
	Add51,
	in_ready_hold,
	stateST_COMP_TRANS,
	mem_used_1,
	in_data_reg_69,
	in_narrow_reg1,
	cp_ready,
	cp_ready1,
	nxt_out_eop,
	out_valid_reg1,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready,
	altera_reset_synchronizer_int_chain_out,
	Decoder1,
	Add2,
	Add21,
	Add22,
	Add23,
	nxt_in_ready1,
	src_valid,
	out_byte_cnt_reg_2,
	cp_ready2,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_6,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	Selector10,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	nxt_out_burstwrap_1,
	nxt_addr_2,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARADDR_0;
input 	h2f_ARADDR_1;
input 	h2f_ARADDR_2;
input 	h2f_ARADDR_3;
input 	h2f_ARBURST_0;
input 	h2f_ARBURST_1;
input 	[128:0] sink0_data;
input 	h2f_ARLEN_0;
input 	Add5;
input 	Add51;
input 	in_ready_hold;
output 	stateST_COMP_TRANS;
input 	mem_used_1;
output 	in_data_reg_69;
output 	in_narrow_reg1;
input 	cp_ready;
input 	cp_ready1;
output 	nxt_out_eop;
output 	out_valid_reg1;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready;
input 	altera_reset_synchronizer_int_chain_out;
input 	Decoder1;
input 	Add2;
input 	Add21;
input 	Add22;
input 	Add23;
output 	nxt_in_ready1;
input 	src_valid;
output 	out_byte_cnt_reg_2;
input 	cp_ready2;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_6;
output 	in_data_reg_105;
output 	in_data_reg_106;
output 	in_data_reg_107;
output 	in_data_reg_108;
output 	in_data_reg_109;
output 	in_data_reg_110;
output 	in_data_reg_111;
output 	in_data_reg_112;
output 	in_data_reg_113;
output 	in_data_reg_114;
output 	in_data_reg_115;
output 	in_data_reg_116;
input 	Selector10;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
input 	nxt_out_burstwrap_1;
input 	nxt_addr_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \align_address_to_size|LessThan0~0_combout ;
wire \align_address_to_size|LessThan0~1_combout ;
wire \nxt_uncomp_subburst_byte_cnt~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt[3]~1_combout ;
wire \nxt_uncomp_subburst_byte_cnt[4]~2_combout ;
wire \Add4~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt[5]~3_combout ;
wire \nxt_uncomp_subburst_byte_cnt[6]~4_combout ;
wire \nxt_uncomp_subburst_byte_cnt[2]~5_combout ;
wire \WideNor1~combout ;
wire \Selector2~1_combout ;
wire \load_next_out_cmd~combout ;
wire \state.ST_UNCOMP_TRANS~q ;
wire \Selector2~0_combout ;
wire \Selector0~0_combout ;
wire \state.ST_IDLE~q ;
wire \Selector1~0_combout ;
wire \Selector1~1_combout ;
wire \NON_PIPELINED_INPUTS.load_next_cmd~0_combout ;
wire \int_bytes_remaining_reg[6]~q ;
wire \d0_int_bytes_remaining[2]~1_combout ;
wire \int_bytes_remaining_reg[2]~q ;
wire \d0_int_bytes_remaining[3]~2_combout ;
wire \int_bytes_remaining_reg[3]~q ;
wire \Add1~1_combout ;
wire \d0_int_bytes_remaining[4]~3_combout ;
wire \int_bytes_remaining_reg[4]~q ;
wire \Add1~0_combout ;
wire \d0_int_bytes_remaining[5]~4_combout ;
wire \int_bytes_remaining_reg[5]~q ;
wire \d0_int_bytes_remaining[6]~0_combout ;
wire \new_burst_reg~0_combout ;
wire \new_burst_reg~q ;
wire \in_bytecount_reg_zero~0_combout ;
wire \in_bytecount_reg_zero~q ;
wire \nxt_out_valid~0_combout ;
wire \nxt_out_valid~1_combout ;
wire \Selector3~0_combout ;
wire \in_burstwrap_reg[3]~q ;
wire \nxt_addr[3]~0_combout ;
wire \nxt_addr[3]~combout ;
wire \int_nxt_addr_reg[3]~q ;
wire \in_size_reg[0]~q ;
wire \in_size_reg[2]~q ;
wire \in_size_reg[1]~q ;
wire \ShiftLeft0~0_combout ;
wire \ShiftLeft0~1_combout ;
wire \int_byte_cnt_narrow_reg[3]~q ;
wire \ShiftLeft0~2_combout ;
wire \int_byte_cnt_narrow_reg[2]~q ;
wire \in_burstwrap_reg[1]~q ;
wire \nxt_addr[1]~combout ;
wire \int_nxt_addr_reg[1]~q ;
wire \ShiftLeft0~3_combout ;
wire \int_byte_cnt_narrow_reg[1]~q ;
wire \int_byte_cnt_narrow_reg[0]~q ;
wire \Add0~13_sumout ;
wire \in_burstwrap_reg[0]~q ;
wire \nxt_addr[0]~combout ;
wire \int_nxt_addr_reg[0]~q ;
wire \d0_int_nxt_addr[0]~2_combout ;
wire \d0_int_nxt_addr[0]~3_combout ;
wire \int_nxt_addr_reg_dly[0]~q ;
wire \Add0~14 ;
wire \Add0~9_sumout ;
wire \d0_int_nxt_addr[1]~4_combout ;
wire \int_nxt_addr_reg_dly[1]~q ;
wire \Add0~10 ;
wire \Add0~6 ;
wire \Add0~1_sumout ;
wire \d0_int_nxt_addr[3]~0_combout ;
wire \in_burstwrap_reg[2]~q ;
wire \nxt_addr[2]~1_combout ;
wire \nxt_addr[2]~combout ;
wire \int_nxt_addr_reg[2]~q ;
wire \Add0~5_sumout ;
wire \d0_int_nxt_addr[2]~1_combout ;


spw_babasu_altera_merlin_address_alignment_2 align_address_to_size(
	.new_burst_reg(\new_burst_reg~q ),
	.src_payload(sink0_data[86]),
	.in_size_reg_0(\in_size_reg[0]~q ),
	.src_payload1(sink0_data[88]),
	.in_size_reg_2(\in_size_reg[2]~q ),
	.src_payload2(sink0_data[87]),
	.in_size_reg_1(\in_size_reg[1]~q ),
	.LessThan0(\align_address_to_size|LessThan0~0_combout ),
	.LessThan01(\align_address_to_size|LessThan0~1_combout ));

dffeas \state.ST_COMP_TRANS (
	.clk(clk_clk),
	.d(\Selector1~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_COMP_TRANS),
	.prn(vcc));
defparam \state.ST_COMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_COMP_TRANS .power_up = "low";

dffeas \in_data_reg[69] (
	.clk(clk_clk),
	.d(sink0_data[69]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_69),
	.prn(vcc));
defparam \in_data_reg[69] .is_wysiwyg = "true";
defparam \in_data_reg[69] .power_up = "low";

dffeas in_narrow_reg(
	.clk(clk_clk),
	.d(Decoder1),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_narrow_reg1),
	.prn(vcc));
defparam in_narrow_reg.is_wysiwyg = "true";
defparam in_narrow_reg.power_up = "low";

cyclonev_lcell_comb \nxt_out_eop~0 (
	.dataa(!in_data_reg_69),
	.datab(!stateST_COMP_TRANS),
	.datac(!\new_burst_reg~q ),
	.datad(!mem_used_1),
	.datae(!cp_ready),
	.dataf(!\in_bytecount_reg_zero~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_out_eop),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_eop~0 .extended_lut = "off";
defparam \nxt_out_eop~0 .lut_mask = 64'h4444474477774777;
defparam \nxt_out_eop~0 .shared_arith = "off";

dffeas out_valid_reg(
	.clk(clk_clk),
	.d(\nxt_out_valid~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_valid_reg1),
	.prn(vcc));
defparam out_valid_reg.is_wysiwyg = "true";
defparam out_valid_reg.power_up = "low";

dffeas \state.ST_UNCOMP_WR_SUBBURST (
	.clk(clk_clk),
	.d(\Selector3~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_UNCOMP_WR_SUBBURST),
	.prn(vcc));
defparam \state.ST_UNCOMP_WR_SUBBURST .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_WR_SUBBURST .power_up = "low";

cyclonev_lcell_comb \nxt_in_ready~0 (
	.dataa(!in_ready_hold),
	.datab(!stateST_COMP_TRANS),
	.datac(!mem_used_1),
	.datad(!cp_ready),
	.datae(!out_valid_reg1),
	.dataf(!\Selector2~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~0 .extended_lut = "off";
defparam \nxt_in_ready~0 .lut_mask = 64'h0000FF3F8888BBBB;
defparam \nxt_in_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_in_ready~1 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!cp_ready1),
	.datac(!nxt_out_eop),
	.datad(!nxt_in_ready),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~1 .extended_lut = "off";
defparam \nxt_in_ready~1 .lut_mask = 64'h00FE00FE00FE00FE;
defparam \nxt_in_ready~1 .shared_arith = "off";

dffeas \out_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[3] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[3]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_3),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[3] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[3] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[2]~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[4] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[4]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_4),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[4] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[4] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[5] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[5]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_5),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[5] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[5] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[6] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[6]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_6),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[6] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[6] .power_up = "low";

dffeas \in_data_reg[105] (
	.clk(clk_clk),
	.d(sink0_data[105]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_105),
	.prn(vcc));
defparam \in_data_reg[105] .is_wysiwyg = "true";
defparam \in_data_reg[105] .power_up = "low";

dffeas \in_data_reg[106] (
	.clk(clk_clk),
	.d(sink0_data[106]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_106),
	.prn(vcc));
defparam \in_data_reg[106] .is_wysiwyg = "true";
defparam \in_data_reg[106] .power_up = "low";

dffeas \in_data_reg[107] (
	.clk(clk_clk),
	.d(sink0_data[107]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_107),
	.prn(vcc));
defparam \in_data_reg[107] .is_wysiwyg = "true";
defparam \in_data_reg[107] .power_up = "low";

dffeas \in_data_reg[108] (
	.clk(clk_clk),
	.d(sink0_data[108]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_108),
	.prn(vcc));
defparam \in_data_reg[108] .is_wysiwyg = "true";
defparam \in_data_reg[108] .power_up = "low";

dffeas \in_data_reg[109] (
	.clk(clk_clk),
	.d(sink0_data[109]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_109),
	.prn(vcc));
defparam \in_data_reg[109] .is_wysiwyg = "true";
defparam \in_data_reg[109] .power_up = "low";

dffeas \in_data_reg[110] (
	.clk(clk_clk),
	.d(sink0_data[110]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_110),
	.prn(vcc));
defparam \in_data_reg[110] .is_wysiwyg = "true";
defparam \in_data_reg[110] .power_up = "low";

dffeas \in_data_reg[111] (
	.clk(clk_clk),
	.d(sink0_data[111]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_111),
	.prn(vcc));
defparam \in_data_reg[111] .is_wysiwyg = "true";
defparam \in_data_reg[111] .power_up = "low";

dffeas \in_data_reg[112] (
	.clk(clk_clk),
	.d(sink0_data[112]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_112),
	.prn(vcc));
defparam \in_data_reg[112] .is_wysiwyg = "true";
defparam \in_data_reg[112] .power_up = "low";

dffeas \in_data_reg[113] (
	.clk(clk_clk),
	.d(sink0_data[113]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_113),
	.prn(vcc));
defparam \in_data_reg[113] .is_wysiwyg = "true";
defparam \in_data_reg[113] .power_up = "low";

dffeas \in_data_reg[114] (
	.clk(clk_clk),
	.d(sink0_data[114]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_114),
	.prn(vcc));
defparam \in_data_reg[114] .is_wysiwyg = "true";
defparam \in_data_reg[114] .power_up = "low";

dffeas \in_data_reg[115] (
	.clk(clk_clk),
	.d(sink0_data[115]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_115),
	.prn(vcc));
defparam \in_data_reg[115] .is_wysiwyg = "true";
defparam \in_data_reg[115] .power_up = "low";

dffeas \in_data_reg[116] (
	.clk(clk_clk),
	.d(sink0_data[116]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_116),
	.prn(vcc));
defparam \in_data_reg[116] .is_wysiwyg = "true";
defparam \in_data_reg[116] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[3] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[3]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_3),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[3] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[2] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[2]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_2),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[2] .power_up = "low";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt~0 (
	.dataa(!cp_ready1),
	.datab(!out_valid_reg1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt~0 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt~0 .lut_mask = 64'h1111111111111111;
defparam \nxt_uncomp_subburst_byte_cnt~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[3]~1 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!out_uncomp_byte_cnt_reg_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[3]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[3]~1 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[3]~1 .lut_mask = 64'h0FE40F4E0FE40F4E;
defparam \nxt_uncomp_subburst_byte_cnt[3]~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[4]~2 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!out_uncomp_byte_cnt_reg_2),
	.dataf(!out_uncomp_byte_cnt_reg_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[4]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[4]~2 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[4]~2 .lut_mask = 64'h00E40044FF4EFFEE;
defparam \nxt_uncomp_subburst_byte_cnt[4]~2 .shared_arith = "off";

cyclonev_lcell_comb \Add4~0 (
	.dataa(!out_uncomp_byte_cnt_reg_3),
	.datab(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datac(!out_uncomp_byte_cnt_reg_2),
	.datad(!out_uncomp_byte_cnt_reg_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add4~0 .extended_lut = "off";
defparam \Add4~0 .lut_mask = 64'h2000200020002000;
defparam \Add4~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[5]~3 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_5),
	.datae(!\Add4~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[5]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[5]~3 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[5]~3 .lut_mask = 64'h04FEAE5404FEAE54;
defparam \nxt_uncomp_subburst_byte_cnt[5]~3 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[6]~4 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_5),
	.datae(!\Add4~0_combout ),
	.dataf(!out_uncomp_byte_cnt_reg_6),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[6]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[6]~4 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[6]~4 .lut_mask = 64'h0404AE04FEFE54FE;
defparam \nxt_uncomp_subburst_byte_cnt[6]~4 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[2]~5 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[2]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[2]~5 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[2]~5 .lut_mask = 64'h0EF40EF40EF40EF4;
defparam \nxt_uncomp_subburst_byte_cnt[2]~5 .shared_arith = "off";

cyclonev_lcell_comb WideNor1(
	.dataa(!\nxt_uncomp_subburst_byte_cnt[3]~1_combout ),
	.datab(!\nxt_uncomp_subburst_byte_cnt[4]~2_combout ),
	.datac(!\nxt_uncomp_subburst_byte_cnt[5]~3_combout ),
	.datad(!\nxt_uncomp_subburst_byte_cnt[6]~4_combout ),
	.datae(!\nxt_uncomp_subburst_byte_cnt[2]~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideNor1.extended_lut = "off";
defparam WideNor1.lut_mask = 64'h8000000080000000;
defparam WideNor1.shared_arith = "off";

cyclonev_lcell_comb \Selector2~1 (
	.dataa(!nxt_out_eop),
	.datab(!\Selector2~0_combout ),
	.datac(!\WideNor1~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~1 .extended_lut = "off";
defparam \Selector2~1 .lut_mask = 64'h0808080808080808;
defparam \Selector2~1 .shared_arith = "off";

cyclonev_lcell_comb load_next_out_cmd(
	.dataa(!mem_used_1),
	.datab(!cp_ready),
	.datac(!out_valid_reg1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\load_next_out_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam load_next_out_cmd.extended_lut = "off";
defparam load_next_out_cmd.lut_mask = 64'hF2F2F2F2F2F2F2F2;
defparam load_next_out_cmd.shared_arith = "off";

dffeas \state.ST_UNCOMP_TRANS (
	.clk(clk_clk),
	.d(\Selector2~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_UNCOMP_TRANS~q ),
	.prn(vcc));
defparam \state.ST_UNCOMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_TRANS .power_up = "low";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'h8888888888888888;
defparam \Selector2~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!in_ready_hold),
	.datab(!nxt_out_eop),
	.datac(!src_valid),
	.datad(!\state.ST_IDLE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'h05CD05CD05CD05CD;
defparam \Selector0~0 .shared_arith = "off";

dffeas \state.ST_IDLE (
	.clk(clk_clk),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_IDLE~q ),
	.prn(vcc));
defparam \state.ST_IDLE .is_wysiwyg = "true";
defparam \state.ST_IDLE .power_up = "low";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!sink0_data[69]),
	.datab(!nxt_out_eop),
	.datac(!\Selector2~0_combout ),
	.datad(!\state.ST_IDLE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'h5510551055105510;
defparam \Selector1~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~1 (
	.dataa(!in_ready_hold),
	.datab(!stateST_COMP_TRANS),
	.datac(!nxt_out_eop),
	.datad(!src_valid),
	.datae(!\Selector1~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~1 .extended_lut = "off";
defparam \Selector1~1 .lut_mask = 64'h3031307530313075;
defparam \Selector1~1 .shared_arith = "off";

cyclonev_lcell_comb \NON_PIPELINED_INPUTS.load_next_cmd~0 (
	.dataa(!in_ready_hold),
	.datab(!nxt_in_ready1),
	.datac(!src_valid),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \NON_PIPELINED_INPUTS.load_next_cmd~0 .extended_lut = "off";
defparam \NON_PIPELINED_INPUTS.load_next_cmd~0 .lut_mask = 64'h0404040404040404;
defparam \NON_PIPELINED_INPUTS.load_next_cmd~0 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[6] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[6]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[6]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[6] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[6] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[2]~1 (
	.dataa(!h2f_ARLEN_0),
	.datab(!sink0_data[69]),
	.datac(!\new_burst_reg~q ),
	.datad(!out_byte_cnt_reg_2),
	.datae(!\int_bytes_remaining_reg[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[2]~1 .extended_lut = "off";
defparam \d0_int_bytes_remaining[2]~1 .lut_mask = 64'h02F2F20202F2F202;
defparam \d0_int_bytes_remaining[2]~1 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[2] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[2]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[2]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[2] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[3]~2 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!Add2),
	.datad(!\int_bytes_remaining_reg[3]~q ),
	.datae(!out_byte_cnt_reg_2),
	.dataf(!\int_bytes_remaining_reg[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[3]~2 .extended_lut = "off";
defparam \d0_int_bytes_remaining[3]~2 .lut_mask = 64'h01CDCD0101CD01CD;
defparam \d0_int_bytes_remaining[3]~2 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[3] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[3]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[3]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[3] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[3] .power_up = "low";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!\int_bytes_remaining_reg[4]~q ),
	.datab(!\int_bytes_remaining_reg[3]~q ),
	.datac(!out_byte_cnt_reg_2),
	.datad(!\int_bytes_remaining_reg[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'hA6AAA6AAA6AAA6AA;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[4]~3 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!Add21),
	.datad(!\Add1~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[4]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[4]~3 .extended_lut = "off";
defparam \d0_int_bytes_remaining[4]~3 .lut_mask = 64'hCD01CD01CD01CD01;
defparam \d0_int_bytes_remaining[4]~3 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[4] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[4]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[4]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[4] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[4] .power_up = "low";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!\int_bytes_remaining_reg[4]~q ),
	.datab(!\int_bytes_remaining_reg[3]~q ),
	.datac(!out_byte_cnt_reg_2),
	.datad(!\int_bytes_remaining_reg[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h0800080008000800;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[5]~4 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!Add22),
	.datad(!\int_bytes_remaining_reg[5]~q ),
	.datae(!\Add1~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[5]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[5]~4 .extended_lut = "off";
defparam \d0_int_bytes_remaining[5]~4 .lut_mask = 64'h01CDCD0101CDCD01;
defparam \d0_int_bytes_remaining[5]~4 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[5] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[5]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[5]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[5] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[5] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[6]~0 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!Add23),
	.datad(!\int_bytes_remaining_reg[6]~q ),
	.datae(!\int_bytes_remaining_reg[5]~q ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[6]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[6]~0 .extended_lut = "off";
defparam \d0_int_bytes_remaining[6]~0 .lut_mask = 64'h01CD01CDCD0101CD;
defparam \d0_int_bytes_remaining[6]~0 .shared_arith = "off";

cyclonev_lcell_comb \new_burst_reg~0 (
	.dataa(!\Selector1~1_combout ),
	.datab(!\d0_int_bytes_remaining[6]~0_combout ),
	.datac(!\d0_int_bytes_remaining[2]~1_combout ),
	.datad(!\d0_int_bytes_remaining[3]~2_combout ),
	.datae(!\d0_int_bytes_remaining[4]~3_combout ),
	.dataf(!\d0_int_bytes_remaining[5]~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\new_burst_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \new_burst_reg~0 .extended_lut = "off";
defparam \new_burst_reg~0 .lut_mask = 64'hAEAAAAAAAAAAAAAA;
defparam \new_burst_reg~0 .shared_arith = "off";

dffeas new_burst_reg(
	.clk(clk_clk),
	.d(\new_burst_reg~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\new_burst_reg~q ),
	.prn(vcc));
defparam new_burst_reg.is_wysiwyg = "true";
defparam new_burst_reg.power_up = "low";

cyclonev_lcell_comb \in_bytecount_reg_zero~0 (
	.dataa(!sink0_data[69]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\in_bytecount_reg_zero~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \in_bytecount_reg_zero~0 .extended_lut = "off";
defparam \in_bytecount_reg_zero~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \in_bytecount_reg_zero~0 .shared_arith = "off";

dffeas in_bytecount_reg_zero(
	.clk(clk_clk),
	.d(\in_bytecount_reg_zero~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_bytecount_reg_zero~q ),
	.prn(vcc));
defparam in_bytecount_reg_zero.is_wysiwyg = "true";
defparam in_bytecount_reg_zero.power_up = "low";

cyclonev_lcell_comb \nxt_out_valid~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!mem_used_1),
	.datac(!\in_bytecount_reg_zero~q ),
	.datad(!cp_ready2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_valid~0 .extended_lut = "off";
defparam \nxt_out_valid~0 .lut_mask = 64'hF0B8F0B8F0B8F0B8;
defparam \nxt_out_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_out_valid~1 (
	.dataa(!in_ready_hold),
	.datab(!stateST_COMP_TRANS),
	.datac(!src_valid),
	.datad(!\nxt_out_valid~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_valid~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_valid~1 .extended_lut = "off";
defparam \nxt_out_valid~1 .lut_mask = 64'h0537053705370537;
defparam \nxt_out_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~0 (
	.dataa(!nxt_out_eop),
	.datab(!\Selector2~0_combout ),
	.datac(!\WideNor1~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'h8080808080808080;
defparam \Selector3~0 .shared_arith = "off";

dffeas \in_burstwrap_reg[3] (
	.clk(clk_clk),
	.d(sink0_data[82]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_burstwrap_reg[3]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[3] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[3] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[3]~0 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!\in_burstwrap_reg[3]~q ),
	.datad(!\d0_int_nxt_addr[3]~0_combout ),
	.datae(!h2f_ARBURST_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[3]~0 .extended_lut = "off";
defparam \nxt_addr[3]~0 .lut_mask = 64'h00F300E200F300E2;
defparam \nxt_addr[3]~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_addr[3] (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!h2f_ARBURST_1),
	.datad(!Add5),
	.datae(!Selector10),
	.dataf(!\nxt_addr[3]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[3] .extended_lut = "off";
defparam \nxt_addr[3] .lut_mask = 64'h00000000FEEEFFEF;
defparam \nxt_addr[3] .shared_arith = "off";

dffeas \int_nxt_addr_reg[3] (
	.clk(clk_clk),
	.d(\nxt_addr[3]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[3]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[3] .power_up = "low";

dffeas \in_size_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[86]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_size_reg[0]~q ),
	.prn(vcc));
defparam \in_size_reg[0] .is_wysiwyg = "true";
defparam \in_size_reg[0] .power_up = "low";

dffeas \in_size_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[88]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_size_reg[2]~q ),
	.prn(vcc));
defparam \in_size_reg[2] .is_wysiwyg = "true";
defparam \in_size_reg[2] .power_up = "low";

dffeas \in_size_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[87]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_size_reg[1]~q ),
	.prn(vcc));
defparam \in_size_reg[1] .is_wysiwyg = "true";
defparam \in_size_reg[1] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[88]),
	.datac(!\in_size_reg[2]~q ),
	.datad(!sink0_data[87]),
	.datae(!\in_size_reg[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~0 .extended_lut = "off";
defparam \ShiftLeft0~0 .lut_mask = 64'h0044A0E40044A0E4;
defparam \ShiftLeft0~0 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~1 .extended_lut = "off";
defparam \ShiftLeft0~1 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~1 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[3] (
	.clk(clk_clk),
	.d(\ShiftLeft0~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[3]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[3] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[3] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~2 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~2 .extended_lut = "off";
defparam \ShiftLeft0~2 .lut_mask = 64'h00E400E400E400E4;
defparam \ShiftLeft0~2 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[2] (
	.clk(clk_clk),
	.d(\ShiftLeft0~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[2]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[2] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[2] .power_up = "low";

dffeas \in_burstwrap_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[80]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_burstwrap_reg[1]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[1] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[1] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[1] (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!\in_burstwrap_reg[1]~q ),
	.datad(!\d0_int_nxt_addr[1]~4_combout ),
	.datae(!nxt_out_burstwrap_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[1] .extended_lut = "off";
defparam \nxt_addr[1] .lut_mask = 64'h00E200F300E200F3;
defparam \nxt_addr[1] .shared_arith = "off";

dffeas \int_nxt_addr_reg[1] (
	.clk(clk_clk),
	.d(\nxt_addr[1]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[1] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\align_address_to_size|LessThan0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~3 .extended_lut = "off";
defparam \ShiftLeft0~3 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~3 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[1] (
	.clk(clk_clk),
	.d(\ShiftLeft0~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[1]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[1] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[1] .power_up = "low";

dffeas \int_byte_cnt_narrow_reg[0] (
	.clk(clk_clk),
	.d(\align_address_to_size|LessThan0~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[0]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[0] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[0] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[0]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \in_burstwrap_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[79]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_burstwrap_reg[0]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[0] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[0] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[0] (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!sink0_data[79]),
	.datad(!\in_burstwrap_reg[0]~q ),
	.datae(!\d0_int_nxt_addr[0]~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[0] .extended_lut = "off";
defparam \nxt_addr[0] .lut_mask = 64'h0000FE320000FE32;
defparam \nxt_addr[0] .shared_arith = "off";

dffeas \int_nxt_addr_reg[0] (
	.clk(clk_clk),
	.d(\nxt_addr[0]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[0] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~2 (
	.dataa(!\Add0~13_sumout ),
	.datab(!\int_nxt_addr_reg[0]~q ),
	.datac(!\in_burstwrap_reg[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~2 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~2 .lut_mask = 64'hC8C8C8C8C8C8C8C8;
defparam \d0_int_nxt_addr[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~3 (
	.dataa(!h2f_ARADDR_0),
	.datab(!sink0_data[69]),
	.datac(!\new_burst_reg~q ),
	.datad(!\align_address_to_size|LessThan0~1_combout ),
	.datae(!\d0_int_nxt_addr[0]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~3 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~3 .lut_mask = 64'hF0F10001F0F10001;
defparam \d0_int_nxt_addr[0]~3 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[0] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[0]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[0] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[1]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[1]~q ),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~4 (
	.dataa(!\int_nxt_addr_reg[1]~q ),
	.datab(!\Add0~9_sumout ),
	.datac(!sink0_data[69]),
	.datad(!Decoder1),
	.datae(!\new_burst_reg~q ),
	.dataf(!h2f_ARADDR_1),
	.datag(!\in_burstwrap_reg[1]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~4 .extended_lut = "on";
defparam \d0_int_nxt_addr[1]~4 .lut_mask = 64'h575700005757000F;
defparam \d0_int_nxt_addr[1]~4 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[1] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[1]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[1] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_2),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[2]~q ),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[3]~q ),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~0 (
	.dataa(!h2f_ARADDR_3),
	.datab(!sink0_data[69]),
	.datac(!\new_burst_reg~q ),
	.datad(!\int_nxt_addr_reg[3]~q ),
	.datae(!\in_burstwrap_reg[3]~q ),
	.dataf(!\Add0~1_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~0 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~0 .lut_mask = 64'h01F101F101F1F1F1;
defparam \d0_int_nxt_addr[3]~0 .shared_arith = "off";

dffeas \in_burstwrap_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[81]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_burstwrap_reg[2]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[2] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[2] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[2]~1 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!\in_burstwrap_reg[2]~q ),
	.datad(!\d0_int_nxt_addr[2]~1_combout ),
	.datae(!h2f_ARBURST_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[2]~1 .extended_lut = "off";
defparam \nxt_addr[2]~1 .lut_mask = 64'h00F300E200F300E2;
defparam \nxt_addr[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_addr[2] (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!h2f_ARBURST_1),
	.datad(!Add51),
	.datae(!\nxt_addr[2]~1_combout ),
	.dataf(!nxt_addr_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[2] .extended_lut = "off";
defparam \nxt_addr[2] .lut_mask = 64'h0000FEEE0000FFEF;
defparam \nxt_addr[2] .shared_arith = "off";

dffeas \int_nxt_addr_reg[2] (
	.clk(clk_clk),
	.d(\nxt_addr[2]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[2]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~1 (
	.dataa(!h2f_ARADDR_2),
	.datab(!sink0_data[69]),
	.datac(!\new_burst_reg~q ),
	.datad(!\int_nxt_addr_reg[2]~q ),
	.datae(!\in_burstwrap_reg[2]~q ),
	.dataf(!\Add0~5_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~1 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~1 .lut_mask = 64'h01F101F101F1F1F1;
defparam \d0_int_nxt_addr[2]~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_address_alignment_2 (
	new_burst_reg,
	src_payload,
	in_size_reg_0,
	src_payload1,
	in_size_reg_2,
	src_payload2,
	in_size_reg_1,
	LessThan0,
	LessThan01)/* synthesis synthesis_greybox=0 */;
input 	new_burst_reg;
input 	src_payload;
input 	in_size_reg_0;
input 	src_payload1;
input 	in_size_reg_2;
input 	src_payload2;
input 	in_size_reg_1;
output 	LessThan0;
output 	LessThan01;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!new_burst_reg),
	.datab(!src_payload1),
	.datac(!in_size_reg_2),
	.datad(!src_payload2),
	.datae(!in_size_reg_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan0),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'hE4A04400E4A04400;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~1 (
	.dataa(!new_burst_reg),
	.datab(!src_payload),
	.datac(!in_size_reg_0),
	.datad(!LessThan0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan01),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~1 .extended_lut = "off";
defparam \LessThan0~1 .lut_mask = 64'h00E400E400E400E4;
defparam \LessThan0~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_burst_adapter_2 (
	h2f_ARADDR_0,
	h2f_ARADDR_1,
	h2f_ARADDR_2,
	h2f_ARADDR_3,
	h2f_ARLEN_0,
	nxt_in_ready,
	in_ready_hold,
	stateST_COMP_TRANS,
	out_valid_reg,
	in_narrow_reg,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	in_data_reg_68,
	cp_ready,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready1,
	saved_grant_1,
	Equal5,
	saved_grant_0,
	altera_reset_synchronizer_int_chain_out,
	in_data_reg_0,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	in_data_reg_1,
	in_data_reg_2,
	in_data_reg_3,
	in_data_reg_4,
	in_data_reg_5,
	in_data_reg_6,
	in_data_reg_7,
	in_data_reg_8,
	Add2,
	Add21,
	Add22,
	Add23,
	Equal51,
	write_cp_data_77,
	write_cp_data_78,
	write_cp_data_75,
	write_cp_data_74,
	write_cp_data_76,
	WideNor0,
	nxt_out_eop,
	src5_valid,
	src_valid,
	cp_ready1,
	in_data_reg_69,
	src_data_87,
	src_data_88,
	src_valid1,
	src_data_35,
	src_data_34,
	src_data_33,
	src_data_32,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_6,
	src_payload_0,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	Selector3,
	Selector10,
	base_address_3,
	Selector4,
	Selector11,
	base_address_2,
	src_payload,
	src_data_82,
	src_data_81,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_data_105,
	src_data_106,
	src_data_107,
	src_data_108,
	src_data_109,
	src_data_110,
	src_data_111,
	src_data_112,
	src_data_113,
	src_data_114,
	src_data_115,
	src_data_116,
	src_data_86,
	Selector5,
	Selector12,
	out_data_1,
	src_data_80,
	out_data_0,
	Selector6,
	Selector13,
	src_data_79,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARADDR_0;
input 	h2f_ARADDR_1;
input 	h2f_ARADDR_2;
input 	h2f_ARADDR_3;
input 	h2f_ARLEN_0;
output 	nxt_in_ready;
input 	in_ready_hold;
output 	stateST_COMP_TRANS;
output 	out_valid_reg;
output 	in_narrow_reg;
output 	in_byteen_reg_3;
output 	in_byteen_reg_2;
output 	in_byteen_reg_1;
output 	in_byteen_reg_0;
output 	in_data_reg_68;
input 	cp_ready;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready1;
input 	saved_grant_1;
input 	Equal5;
input 	saved_grant_0;
input 	altera_reset_synchronizer_int_chain_out;
output 	in_data_reg_0;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
output 	in_data_reg_1;
output 	in_data_reg_2;
output 	in_data_reg_3;
output 	in_data_reg_4;
output 	in_data_reg_5;
output 	in_data_reg_6;
output 	in_data_reg_7;
output 	in_data_reg_8;
input 	Add2;
input 	Add21;
input 	Add22;
input 	Add23;
input 	Equal51;
input 	write_cp_data_77;
input 	write_cp_data_78;
input 	write_cp_data_75;
input 	write_cp_data_74;
input 	write_cp_data_76;
input 	WideNor0;
output 	nxt_out_eop;
input 	src5_valid;
input 	src_valid;
input 	cp_ready1;
output 	in_data_reg_69;
input 	src_data_87;
input 	src_data_88;
input 	src_valid1;
input 	src_data_35;
input 	src_data_34;
input 	src_data_33;
input 	src_data_32;
output 	out_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_6;
input 	src_payload_0;
output 	in_data_reg_105;
output 	in_data_reg_106;
output 	in_data_reg_107;
output 	in_data_reg_108;
output 	in_data_reg_109;
output 	in_data_reg_110;
output 	in_data_reg_111;
output 	in_data_reg_112;
output 	in_data_reg_113;
output 	in_data_reg_114;
output 	in_data_reg_115;
output 	in_data_reg_116;
input 	Selector3;
input 	Selector10;
input 	base_address_3;
input 	Selector4;
input 	Selector11;
input 	base_address_2;
input 	src_payload;
input 	src_data_82;
input 	src_data_81;
input 	src_payload1;
input 	src_payload2;
input 	src_payload3;
input 	src_payload4;
input 	src_payload5;
input 	src_payload6;
input 	src_payload7;
input 	src_payload8;
input 	src_data_105;
input 	src_data_106;
input 	src_data_107;
input 	src_data_108;
input 	src_data_109;
input 	src_data_110;
input 	src_data_111;
input 	src_data_112;
input 	src_data_113;
input 	src_data_114;
input 	src_data_115;
input 	src_data_116;
input 	src_data_86;
input 	Selector5;
input 	Selector12;
input 	out_data_1;
input 	src_data_80;
input 	out_data_0;
input 	Selector6;
input 	Selector13;
input 	src_data_79;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



spw_babasu_altera_merlin_burst_adapter_13_1_2 \altera_merlin_burst_adapter_13_1.burst_adapter (
	.h2f_ARADDR_0(h2f_ARADDR_0),
	.h2f_ARADDR_1(h2f_ARADDR_1),
	.h2f_ARADDR_2(h2f_ARADDR_2),
	.h2f_ARADDR_3(h2f_ARADDR_3),
	.h2f_ARLEN_0(h2f_ARLEN_0),
	.nxt_in_ready(nxt_in_ready),
	.in_ready_hold(in_ready_hold),
	.stateST_COMP_TRANS(stateST_COMP_TRANS),
	.out_valid_reg1(out_valid_reg),
	.in_narrow_reg1(in_narrow_reg),
	.in_byteen_reg_3(in_byteen_reg_3),
	.in_byteen_reg_2(in_byteen_reg_2),
	.in_byteen_reg_1(in_byteen_reg_1),
	.in_byteen_reg_0(in_byteen_reg_0),
	.in_data_reg_68(in_data_reg_68),
	.cp_ready(cp_ready),
	.stateST_UNCOMP_WR_SUBBURST(stateST_UNCOMP_WR_SUBBURST),
	.nxt_in_ready1(nxt_in_ready1),
	.sink0_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_116,src_data_115,src_data_114,src_data_113,src_data_112,src_data_111,src_data_110,src_data_109,src_data_108,src_data_107,src_data_106,src_data_105,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_88,src_data_87,
src_data_86,gnd,gnd,gnd,src_data_82,src_data_81,src_data_80,src_data_79,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,saved_grant_1,saved_grant_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_35,src_data_34,src_data_33,
src_data_32,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_payload8,src_payload7,src_payload6,src_payload5,src_payload4,src_payload3,src_payload2,src_payload1,src_payload}),
	.Equal5(Equal5),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.in_data_reg_0(in_data_reg_0),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_3),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_2),
	.in_data_reg_1(in_data_reg_1),
	.in_data_reg_2(in_data_reg_2),
	.in_data_reg_3(in_data_reg_3),
	.in_data_reg_4(in_data_reg_4),
	.in_data_reg_5(in_data_reg_5),
	.in_data_reg_6(in_data_reg_6),
	.in_data_reg_7(in_data_reg_7),
	.in_data_reg_8(in_data_reg_8),
	.Add2(Add2),
	.Add21(Add21),
	.Add22(Add22),
	.Add23(Add23),
	.Equal51(Equal51),
	.write_cp_data_77(write_cp_data_77),
	.write_cp_data_78(write_cp_data_78),
	.write_cp_data_75(write_cp_data_75),
	.write_cp_data_74(write_cp_data_74),
	.write_cp_data_76(write_cp_data_76),
	.WideNor0(WideNor0),
	.nxt_out_eop(nxt_out_eop),
	.src5_valid(src5_valid),
	.src_valid(src_valid),
	.cp_ready1(cp_ready1),
	.in_data_reg_69(in_data_reg_69),
	.src_valid1(src_valid1),
	.out_byte_cnt_reg_2(out_byte_cnt_reg_2),
	.out_uncomp_byte_cnt_reg_3(out_uncomp_byte_cnt_reg_3),
	.out_uncomp_byte_cnt_reg_2(out_uncomp_byte_cnt_reg_2),
	.out_uncomp_byte_cnt_reg_4(out_uncomp_byte_cnt_reg_4),
	.out_uncomp_byte_cnt_reg_5(out_uncomp_byte_cnt_reg_5),
	.out_uncomp_byte_cnt_reg_6(out_uncomp_byte_cnt_reg_6),
	.sink0_endofpacket(src_payload_0),
	.in_data_reg_105(in_data_reg_105),
	.in_data_reg_106(in_data_reg_106),
	.in_data_reg_107(in_data_reg_107),
	.in_data_reg_108(in_data_reg_108),
	.in_data_reg_109(in_data_reg_109),
	.in_data_reg_110(in_data_reg_110),
	.in_data_reg_111(in_data_reg_111),
	.in_data_reg_112(in_data_reg_112),
	.in_data_reg_113(in_data_reg_113),
	.in_data_reg_114(in_data_reg_114),
	.in_data_reg_115(in_data_reg_115),
	.in_data_reg_116(in_data_reg_116),
	.Selector3(Selector3),
	.Selector10(Selector10),
	.base_address_3(base_address_3),
	.Selector4(Selector4),
	.Selector11(Selector11),
	.base_address_2(base_address_2),
	.Selector5(Selector5),
	.Selector12(Selector12),
	.out_data_1(out_data_1),
	.out_data_0(out_data_0),
	.Selector6(Selector6),
	.Selector13(Selector13),
	.clk_clk(clk_clk));

endmodule

module spw_babasu_altera_merlin_burst_adapter_13_1_2 (
	h2f_ARADDR_0,
	h2f_ARADDR_1,
	h2f_ARADDR_2,
	h2f_ARADDR_3,
	h2f_ARLEN_0,
	nxt_in_ready,
	in_ready_hold,
	stateST_COMP_TRANS,
	out_valid_reg1,
	in_narrow_reg1,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	in_data_reg_68,
	cp_ready,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready1,
	sink0_data,
	Equal5,
	altera_reset_synchronizer_int_chain_out,
	in_data_reg_0,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	in_data_reg_1,
	in_data_reg_2,
	in_data_reg_3,
	in_data_reg_4,
	in_data_reg_5,
	in_data_reg_6,
	in_data_reg_7,
	in_data_reg_8,
	Add2,
	Add21,
	Add22,
	Add23,
	Equal51,
	write_cp_data_77,
	write_cp_data_78,
	write_cp_data_75,
	write_cp_data_74,
	write_cp_data_76,
	WideNor0,
	nxt_out_eop,
	src5_valid,
	src_valid,
	cp_ready1,
	in_data_reg_69,
	src_valid1,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_6,
	sink0_endofpacket,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	Selector3,
	Selector10,
	base_address_3,
	Selector4,
	Selector11,
	base_address_2,
	Selector5,
	Selector12,
	out_data_1,
	out_data_0,
	Selector6,
	Selector13,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARADDR_0;
input 	h2f_ARADDR_1;
input 	h2f_ARADDR_2;
input 	h2f_ARADDR_3;
input 	h2f_ARLEN_0;
output 	nxt_in_ready;
input 	in_ready_hold;
output 	stateST_COMP_TRANS;
output 	out_valid_reg1;
output 	in_narrow_reg1;
output 	in_byteen_reg_3;
output 	in_byteen_reg_2;
output 	in_byteen_reg_1;
output 	in_byteen_reg_0;
output 	in_data_reg_68;
input 	cp_ready;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready1;
input 	[128:0] sink0_data;
input 	Equal5;
input 	altera_reset_synchronizer_int_chain_out;
output 	in_data_reg_0;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
output 	in_data_reg_1;
output 	in_data_reg_2;
output 	in_data_reg_3;
output 	in_data_reg_4;
output 	in_data_reg_5;
output 	in_data_reg_6;
output 	in_data_reg_7;
output 	in_data_reg_8;
input 	Add2;
input 	Add21;
input 	Add22;
input 	Add23;
input 	Equal51;
input 	write_cp_data_77;
input 	write_cp_data_78;
input 	write_cp_data_75;
input 	write_cp_data_74;
input 	write_cp_data_76;
input 	WideNor0;
output 	nxt_out_eop;
input 	src5_valid;
input 	src_valid;
input 	cp_ready1;
output 	in_data_reg_69;
input 	src_valid1;
output 	out_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_6;
input 	sink0_endofpacket;
output 	in_data_reg_105;
output 	in_data_reg_106;
output 	in_data_reg_107;
output 	in_data_reg_108;
output 	in_data_reg_109;
output 	in_data_reg_110;
output 	in_data_reg_111;
output 	in_data_reg_112;
output 	in_data_reg_113;
output 	in_data_reg_114;
output 	in_data_reg_115;
output 	in_data_reg_116;
input 	Selector3;
input 	Selector10;
input 	base_address_3;
input 	Selector4;
input 	Selector11;
input 	base_address_2;
input 	Selector5;
input 	Selector12;
input 	out_data_1;
input 	out_data_0;
input 	Selector6;
input 	Selector13;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \align_address_to_size|LessThan0~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt[3]~1_combout ;
wire \nxt_uncomp_subburst_byte_cnt[4]~2_combout ;
wire \Add4~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt[5]~3_combout ;
wire \nxt_uncomp_subburst_byte_cnt[2]~4_combout ;
wire \nxt_uncomp_subburst_byte_cnt[6]~5_combout ;
wire \WideOr0~combout ;
wire \in_valid~combout ;
wire \Selector0~0_combout ;
wire \load_next_out_cmd~combout ;
wire \state.ST_IDLE~q ;
wire \Selector2~0_combout ;
wire \Selector2~1_combout ;
wire \Selector2~2_combout ;
wire \state.ST_UNCOMP_TRANS~q ;
wire \Selector1~0_combout ;
wire \Selector1~1_combout ;
wire \int_bytes_remaining_reg[3]~q ;
wire \d0_int_bytes_remaining[2]~2_combout ;
wire \d0_int_bytes_remaining[2]~3_combout ;
wire \int_bytes_remaining_reg[2]~q ;
wire \d0_int_bytes_remaining[3]~0_combout ;
wire \d0_int_bytes_remaining[3]~1_combout ;
wire \int_bytes_remaining_reg[6]~q ;
wire \Add1~1_combout ;
wire \d0_int_bytes_remaining[4]~8_combout ;
wire \int_bytes_remaining_reg[4]~q ;
wire \Add1~0_combout ;
wire \d0_int_bytes_remaining[5]~6_combout ;
wire \d0_int_bytes_remaining[5]~7_combout ;
wire \int_bytes_remaining_reg[5]~q ;
wire \d0_int_bytes_remaining[6]~4_combout ;
wire \d0_int_bytes_remaining[6]~5_combout ;
wire \new_burst_reg~0_combout ;
wire \new_burst_reg~q ;
wire \WideNor0~0_combout ;
wire \NON_PIPELINED_INPUTS.load_next_cmd~combout ;
wire \in_bytecount_reg_zero~q ;
wire \nxt_out_valid~0_combout ;
wire \LessThan0~0_combout ;
wire \Selector3~0_combout ;
wire \in_size_reg[0]~q ;
wire \in_size_reg[1]~q ;
wire \in_size_reg[2]~q ;
wire \ShiftLeft0~0_combout ;
wire \ShiftLeft0~1_combout ;
wire \int_byte_cnt_narrow_reg[3]~q ;
wire \ShiftLeft0~2_combout ;
wire \int_byte_cnt_narrow_reg[2]~q ;
wire \ShiftLeft0~3_combout ;
wire \ShiftLeft0~4_combout ;
wire \int_byte_cnt_narrow_reg[1]~q ;
wire \int_byte_cnt_narrow_reg[0]~q ;
wire \Add0~13_sumout ;
wire \d0_int_nxt_addr[0]~3_combout ;
wire \in_burstwrap_reg[0]~q ;
wire \nxt_addr[0]~0_combout ;
wire \int_nxt_addr_reg[0]~q ;
wire \d0_int_nxt_addr[0]~4_combout ;
wire \int_nxt_addr_reg_dly[0]~q ;
wire \Add0~14 ;
wire \Add0~9_sumout ;
wire \in_burstwrap_reg[1]~q ;
wire \nxt_addr[1]~4_combout ;
wire \int_nxt_addr_reg[1]~q ;
wire \d0_int_nxt_addr[1]~7_combout ;
wire \d0_int_nxt_addr[1]~2_combout ;
wire \int_nxt_addr_reg_dly[1]~q ;
wire \Add0~10 ;
wire \Add0~6 ;
wire \Add0~1_sumout ;
wire \in_burstwrap_reg[3]~q ;
wire \nxt_addr[3]~12_combout ;
wire \int_nxt_addr_reg[3]~q ;
wire \d0_int_nxt_addr[3]~5_combout ;
wire \d0_int_nxt_addr[3]~0_combout ;
wire \Add0~5_sumout ;
wire \in_burstwrap_reg[2]~q ;
wire \nxt_addr[2]~8_combout ;
wire \int_nxt_addr_reg[2]~q ;
wire \d0_int_nxt_addr[2]~6_combout ;
wire \d0_int_nxt_addr[2]~1_combout ;
wire \in_eop_reg~q ;


spw_babasu_altera_merlin_address_alignment_3 align_address_to_size(
	.new_burst_reg(\new_burst_reg~q ),
	.src_data_86(sink0_data[86]),
	.in_size_reg_0(\in_size_reg[0]~q ),
	.ShiftLeft0(\ShiftLeft0~3_combout ),
	.LessThan0(\align_address_to_size|LessThan0~0_combout ));

cyclonev_lcell_comb \nxt_in_ready~1 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!in_ready_hold),
	.datac(!out_valid_reg1),
	.datad(!cp_ready),
	.datae(!stateST_COMP_TRANS),
	.dataf(!\new_burst_reg~q ),
	.datag(!stateST_UNCOMP_WR_SUBBURST),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~1 .extended_lut = "on";
defparam \nxt_in_ready~1 .lut_mask = 64'h2020F0F02020F0FF;
defparam \nxt_in_ready~1 .shared_arith = "off";

dffeas \state.ST_COMP_TRANS (
	.clk(clk_clk),
	.d(\Selector1~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_COMP_TRANS),
	.prn(vcc));
defparam \state.ST_COMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_COMP_TRANS .power_up = "low";

dffeas out_valid_reg(
	.clk(clk_clk),
	.d(\nxt_out_valid~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_valid_reg1),
	.prn(vcc));
defparam out_valid_reg.is_wysiwyg = "true";
defparam out_valid_reg.power_up = "low";

dffeas in_narrow_reg(
	.clk(clk_clk),
	.d(\LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_narrow_reg1),
	.prn(vcc));
defparam in_narrow_reg.is_wysiwyg = "true";
defparam in_narrow_reg.power_up = "low";

dffeas \in_byteen_reg[3] (
	.clk(clk_clk),
	.d(sink0_data[35]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_3),
	.prn(vcc));
defparam \in_byteen_reg[3] .is_wysiwyg = "true";
defparam \in_byteen_reg[3] .power_up = "low";

dffeas \in_byteen_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[34]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_2),
	.prn(vcc));
defparam \in_byteen_reg[2] .is_wysiwyg = "true";
defparam \in_byteen_reg[2] .power_up = "low";

dffeas \in_byteen_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[33]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_1),
	.prn(vcc));
defparam \in_byteen_reg[1] .is_wysiwyg = "true";
defparam \in_byteen_reg[1] .power_up = "low";

dffeas \in_byteen_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[32]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_0),
	.prn(vcc));
defparam \in_byteen_reg[0] .is_wysiwyg = "true";
defparam \in_byteen_reg[0] .power_up = "low";

dffeas \in_data_reg[68] (
	.clk(clk_clk),
	.d(sink0_data[68]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_68),
	.prn(vcc));
defparam \in_data_reg[68] .is_wysiwyg = "true";
defparam \in_data_reg[68] .power_up = "low";

dffeas \state.ST_UNCOMP_WR_SUBBURST (
	.clk(clk_clk),
	.d(\Selector3~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_UNCOMP_WR_SUBBURST),
	.prn(vcc));
defparam \state.ST_UNCOMP_WR_SUBBURST .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_WR_SUBBURST .power_up = "low";

cyclonev_lcell_comb \nxt_in_ready~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!out_valid_reg1),
	.datac(!cp_ready),
	.datad(!\state.ST_UNCOMP_TRANS~q ),
	.datae(!stateST_UNCOMP_WR_SUBBURST),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~0 .extended_lut = "off";
defparam \nxt_in_ready~0 .lut_mask = 64'h008A8A8A008A8A8A;
defparam \nxt_in_ready~0 .shared_arith = "off";

dffeas \in_data_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[0]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_0),
	.prn(vcc));
defparam \in_data_reg[0] .is_wysiwyg = "true";
defparam \in_data_reg[0] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[3] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[3]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_3),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[3] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[2] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[2]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_2),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[2] .power_up = "low";

dffeas \in_data_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[1]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_1),
	.prn(vcc));
defparam \in_data_reg[1] .is_wysiwyg = "true";
defparam \in_data_reg[1] .power_up = "low";

dffeas \in_data_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[2]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_2),
	.prn(vcc));
defparam \in_data_reg[2] .is_wysiwyg = "true";
defparam \in_data_reg[2] .power_up = "low";

dffeas \in_data_reg[3] (
	.clk(clk_clk),
	.d(sink0_data[3]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_3),
	.prn(vcc));
defparam \in_data_reg[3] .is_wysiwyg = "true";
defparam \in_data_reg[3] .power_up = "low";

dffeas \in_data_reg[4] (
	.clk(clk_clk),
	.d(sink0_data[4]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_4),
	.prn(vcc));
defparam \in_data_reg[4] .is_wysiwyg = "true";
defparam \in_data_reg[4] .power_up = "low";

dffeas \in_data_reg[5] (
	.clk(clk_clk),
	.d(sink0_data[5]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_5),
	.prn(vcc));
defparam \in_data_reg[5] .is_wysiwyg = "true";
defparam \in_data_reg[5] .power_up = "low";

dffeas \in_data_reg[6] (
	.clk(clk_clk),
	.d(sink0_data[6]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_6),
	.prn(vcc));
defparam \in_data_reg[6] .is_wysiwyg = "true";
defparam \in_data_reg[6] .power_up = "low";

dffeas \in_data_reg[7] (
	.clk(clk_clk),
	.d(sink0_data[7]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_7),
	.prn(vcc));
defparam \in_data_reg[7] .is_wysiwyg = "true";
defparam \in_data_reg[7] .power_up = "low";

dffeas \in_data_reg[8] (
	.clk(clk_clk),
	.d(sink0_data[8]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_8),
	.prn(vcc));
defparam \in_data_reg[8] .is_wysiwyg = "true";
defparam \in_data_reg[8] .power_up = "low";

cyclonev_lcell_comb \nxt_out_eop~0 (
	.dataa(!\in_eop_reg~q ),
	.datab(!stateST_COMP_TRANS),
	.datac(!\new_burst_reg~q ),
	.datad(!cp_ready),
	.datae(!\in_bytecount_reg_zero~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_out_eop),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_eop~0 .extended_lut = "off";
defparam \nxt_out_eop~0 .lut_mask = 64'h4447774744477747;
defparam \nxt_out_eop~0 .shared_arith = "off";

dffeas \in_data_reg[69] (
	.clk(clk_clk),
	.d(sink0_data[69]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_69),
	.prn(vcc));
defparam \in_data_reg[69] .is_wysiwyg = "true";
defparam \in_data_reg[69] .power_up = "low";

dffeas \out_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[3] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[3]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_3),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[3] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[3] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[2]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[4] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[4]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_4),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[4] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[4] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[5] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[5]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_5),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[5] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[5] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[6] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[6]~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_6),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[6] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[6] .power_up = "low";

dffeas \in_data_reg[105] (
	.clk(clk_clk),
	.d(sink0_data[105]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_105),
	.prn(vcc));
defparam \in_data_reg[105] .is_wysiwyg = "true";
defparam \in_data_reg[105] .power_up = "low";

dffeas \in_data_reg[106] (
	.clk(clk_clk),
	.d(sink0_data[106]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_106),
	.prn(vcc));
defparam \in_data_reg[106] .is_wysiwyg = "true";
defparam \in_data_reg[106] .power_up = "low";

dffeas \in_data_reg[107] (
	.clk(clk_clk),
	.d(sink0_data[107]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_107),
	.prn(vcc));
defparam \in_data_reg[107] .is_wysiwyg = "true";
defparam \in_data_reg[107] .power_up = "low";

dffeas \in_data_reg[108] (
	.clk(clk_clk),
	.d(sink0_data[108]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_108),
	.prn(vcc));
defparam \in_data_reg[108] .is_wysiwyg = "true";
defparam \in_data_reg[108] .power_up = "low";

dffeas \in_data_reg[109] (
	.clk(clk_clk),
	.d(sink0_data[109]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_109),
	.prn(vcc));
defparam \in_data_reg[109] .is_wysiwyg = "true";
defparam \in_data_reg[109] .power_up = "low";

dffeas \in_data_reg[110] (
	.clk(clk_clk),
	.d(sink0_data[110]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_110),
	.prn(vcc));
defparam \in_data_reg[110] .is_wysiwyg = "true";
defparam \in_data_reg[110] .power_up = "low";

dffeas \in_data_reg[111] (
	.clk(clk_clk),
	.d(sink0_data[111]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_111),
	.prn(vcc));
defparam \in_data_reg[111] .is_wysiwyg = "true";
defparam \in_data_reg[111] .power_up = "low";

dffeas \in_data_reg[112] (
	.clk(clk_clk),
	.d(sink0_data[112]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_112),
	.prn(vcc));
defparam \in_data_reg[112] .is_wysiwyg = "true";
defparam \in_data_reg[112] .power_up = "low";

dffeas \in_data_reg[113] (
	.clk(clk_clk),
	.d(sink0_data[113]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_113),
	.prn(vcc));
defparam \in_data_reg[113] .is_wysiwyg = "true";
defparam \in_data_reg[113] .power_up = "low";

dffeas \in_data_reg[114] (
	.clk(clk_clk),
	.d(sink0_data[114]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_114),
	.prn(vcc));
defparam \in_data_reg[114] .is_wysiwyg = "true";
defparam \in_data_reg[114] .power_up = "low";

dffeas \in_data_reg[115] (
	.clk(clk_clk),
	.d(sink0_data[115]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_115),
	.prn(vcc));
defparam \in_data_reg[115] .is_wysiwyg = "true";
defparam \in_data_reg[115] .power_up = "low";

dffeas \in_data_reg[116] (
	.clk(clk_clk),
	.d(sink0_data[116]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_116),
	.prn(vcc));
defparam \in_data_reg[116] .is_wysiwyg = "true";
defparam \in_data_reg[116] .power_up = "low";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt~0 (
	.dataa(!out_valid_reg1),
	.datab(!cp_ready),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt~0 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt~0 .lut_mask = 64'h1111111111111111;
defparam \nxt_uncomp_subburst_byte_cnt~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[3]~1 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!out_uncomp_byte_cnt_reg_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[3]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[3]~1 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[3]~1 .lut_mask = 64'h0FE40F4E0FE40F4E;
defparam \nxt_uncomp_subburst_byte_cnt[3]~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[4]~2 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!out_uncomp_byte_cnt_reg_2),
	.dataf(!out_uncomp_byte_cnt_reg_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[4]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[4]~2 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[4]~2 .lut_mask = 64'h00E40044FF4EFFEE;
defparam \nxt_uncomp_subburst_byte_cnt[4]~2 .shared_arith = "off";

cyclonev_lcell_comb \Add4~0 (
	.dataa(!out_uncomp_byte_cnt_reg_3),
	.datab(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datac(!out_uncomp_byte_cnt_reg_2),
	.datad(!out_uncomp_byte_cnt_reg_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add4~0 .extended_lut = "off";
defparam \Add4~0 .lut_mask = 64'h2000200020002000;
defparam \Add4~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[5]~3 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_5),
	.datae(!\Add4~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[5]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[5]~3 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[5]~3 .lut_mask = 64'h04FEAE5404FEAE54;
defparam \nxt_uncomp_subburst_byte_cnt[5]~3 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[2]~4 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[2]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[2]~4 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[2]~4 .lut_mask = 64'h0EF40EF40EF40EF4;
defparam \nxt_uncomp_subburst_byte_cnt[2]~4 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[6]~5 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_5),
	.datae(!\Add4~0_combout ),
	.dataf(!out_uncomp_byte_cnt_reg_6),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[6]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[6]~5 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[6]~5 .lut_mask = 64'h0404AE04FEFE54FE;
defparam \nxt_uncomp_subburst_byte_cnt[6]~5 .shared_arith = "off";

cyclonev_lcell_comb WideOr0(
	.dataa(!\nxt_uncomp_subburst_byte_cnt[3]~1_combout ),
	.datab(!\nxt_uncomp_subburst_byte_cnt[4]~2_combout ),
	.datac(!\nxt_uncomp_subburst_byte_cnt[5]~3_combout ),
	.datad(!\nxt_uncomp_subburst_byte_cnt[2]~4_combout ),
	.datae(!\nxt_uncomp_subburst_byte_cnt[6]~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr0.extended_lut = "off";
defparam WideOr0.lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam WideOr0.shared_arith = "off";

cyclonev_lcell_comb in_valid(
	.dataa(!in_ready_hold),
	.datab(!Equal51),
	.datac(!Equal5),
	.datad(!sink0_data[68]),
	.datae(!src5_valid),
	.dataf(!src_valid),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\in_valid~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam in_valid.extended_lut = "off";
defparam in_valid.lut_mask = 64'h0000000155555555;
defparam in_valid.shared_arith = "off";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!sink0_data[69]),
	.datab(!nxt_out_eop),
	.datac(!sink0_data[68]),
	.datad(!\in_valid~combout ),
	.datae(!\state.ST_IDLE~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'h005FCCFF005FCCFF;
defparam \Selector0~0 .shared_arith = "off";

cyclonev_lcell_comb load_next_out_cmd(
	.dataa(!out_valid_reg1),
	.datab(!cp_ready),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\load_next_out_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam load_next_out_cmd.extended_lut = "off";
defparam load_next_out_cmd.lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam load_next_out_cmd.shared_arith = "off";

dffeas \state.ST_IDLE (
	.clk(clk_clk),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_IDLE~q ),
	.prn(vcc));
defparam \state.ST_IDLE .is_wysiwyg = "true";
defparam \state.ST_IDLE .power_up = "low";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!nxt_out_eop),
	.datac(!stateST_UNCOMP_WR_SUBBURST),
	.datad(!\state.ST_IDLE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'h00EC00EC00EC00EC;
defparam \Selector2~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~1 (
	.dataa(!in_ready_hold),
	.datab(!Equal51),
	.datac(!Equal5),
	.datad(!sink0_data[68]),
	.datae(!src5_valid),
	.dataf(!\Selector2~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~1 .extended_lut = "off";
defparam \Selector2~1 .lut_mask = 64'h0000000100000000;
defparam \Selector2~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~2 (
	.dataa(!\WideOr0~combout ),
	.datab(!\Selector2~1_combout ),
	.datac(!\in_valid~combout ),
	.datad(!nxt_out_eop),
	.datae(!\state.ST_UNCOMP_TRANS~q ),
	.dataf(!sink0_data[69]),
	.datag(!stateST_UNCOMP_WR_SUBBURST),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~2 .extended_lut = "on";
defparam \Selector2~2 .lut_mask = 64'h3B33BB3F0A00AA00;
defparam \Selector2~2 .shared_arith = "off";

dffeas \state.ST_UNCOMP_TRANS (
	.clk(clk_clk),
	.d(\Selector2~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_UNCOMP_TRANS~q ),
	.prn(vcc));
defparam \state.ST_UNCOMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_TRANS .power_up = "low";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!nxt_out_eop),
	.datac(!\state.ST_UNCOMP_TRANS~q ),
	.datad(!stateST_UNCOMP_WR_SUBBURST),
	.datae(!\state.ST_IDLE~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'h0000A8880000A888;
defparam \Selector1~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~1 (
	.dataa(!sink0_data[69]),
	.datab(!stateST_COMP_TRANS),
	.datac(!nxt_out_eop),
	.datad(!sink0_data[68]),
	.datae(!\in_valid~combout ),
	.dataf(!\Selector1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~1 .extended_lut = "off";
defparam \Selector1~1 .lut_mask = 64'h3030777530303330;
defparam \Selector1~1 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[3] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[3]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[3]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[3] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[3] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[2]~2 (
	.dataa(!h2f_ARLEN_0),
	.datab(!sink0_data[69]),
	.datac(!sink0_data[68]),
	.datad(!write_cp_data_74),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[2]~2 .extended_lut = "off";
defparam \d0_int_bytes_remaining[2]~2 .lut_mask = 64'h2F222F222F222F22;
defparam \d0_int_bytes_remaining[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[2]~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\int_bytes_remaining_reg[2]~q ),
	.datad(!\d0_int_bytes_remaining[2]~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[2]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[2]~3 .extended_lut = "off";
defparam \d0_int_bytes_remaining[2]~3 .lut_mask = 64'h287D287D287D287D;
defparam \d0_int_bytes_remaining[2]~3 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[2] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[2]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[2]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[2] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[3]~0 (
	.dataa(!sink0_data[69]),
	.datab(!sink0_data[68]),
	.datac(!write_cp_data_75),
	.datad(!Add2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[3]~0 .extended_lut = "off";
defparam \d0_int_bytes_remaining[3]~0 .lut_mask = 64'h0357035703570357;
defparam \d0_int_bytes_remaining[3]~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[3]~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\int_bytes_remaining_reg[3]~q ),
	.datac(!out_byte_cnt_reg_2),
	.datad(!\int_bytes_remaining_reg[2]~q ),
	.datae(!\d0_int_bytes_remaining[3]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[3]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[3]~1 .extended_lut = "off";
defparam \d0_int_bytes_remaining[3]~1 .lut_mask = 64'h28227D7728227D77;
defparam \d0_int_bytes_remaining[3]~1 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[6] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[6]~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[6]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[6] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[6] .power_up = "low";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!\int_bytes_remaining_reg[3]~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\int_bytes_remaining_reg[2]~q ),
	.datad(!\int_bytes_remaining_reg[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'hDF20DF20DF20DF20;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[4]~8 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!sink0_data[68]),
	.datad(!write_cp_data_76),
	.datae(!Add21),
	.dataf(!\Add1~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[4]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[4]~8 .extended_lut = "off";
defparam \d0_int_bytes_remaining[4]~8 .lut_mask = 64'hCCCFDDDF00031113;
defparam \d0_int_bytes_remaining[4]~8 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[4] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[4]~8_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[4]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[4] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[4] .power_up = "low";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!\int_bytes_remaining_reg[3]~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\int_bytes_remaining_reg[2]~q ),
	.datad(!\int_bytes_remaining_reg[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h2000200020002000;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[5]~6 (
	.dataa(!sink0_data[69]),
	.datab(!sink0_data[68]),
	.datac(!write_cp_data_77),
	.datad(!Add22),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[5]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[5]~6 .extended_lut = "off";
defparam \d0_int_bytes_remaining[5]~6 .lut_mask = 64'h0357035703570357;
defparam \d0_int_bytes_remaining[5]~6 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[5]~7 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\int_bytes_remaining_reg[5]~q ),
	.datac(!\Add1~0_combout ),
	.datad(!\d0_int_bytes_remaining[5]~6_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[5]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[5]~7 .extended_lut = "off";
defparam \d0_int_bytes_remaining[5]~7 .lut_mask = 64'h287D287D287D287D;
defparam \d0_int_bytes_remaining[5]~7 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[5] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[5]~7_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[5]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[5] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[5] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[6]~4 (
	.dataa(!sink0_data[69]),
	.datab(!sink0_data[68]),
	.datac(!write_cp_data_78),
	.datad(!Add23),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[6]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[6]~4 .extended_lut = "off";
defparam \d0_int_bytes_remaining[6]~4 .lut_mask = 64'h0357035703570357;
defparam \d0_int_bytes_remaining[6]~4 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[6]~5 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\int_bytes_remaining_reg[6]~q ),
	.datac(!\int_bytes_remaining_reg[5]~q ),
	.datad(!\Add1~0_combout ),
	.datae(!\d0_int_bytes_remaining[6]~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[6]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[6]~5 .extended_lut = "off";
defparam \d0_int_bytes_remaining[6]~5 .lut_mask = 64'h228277D7228277D7;
defparam \d0_int_bytes_remaining[6]~5 .shared_arith = "off";

cyclonev_lcell_comb \new_burst_reg~0 (
	.dataa(!\Selector1~1_combout ),
	.datab(!\d0_int_bytes_remaining[3]~1_combout ),
	.datac(!\d0_int_bytes_remaining[2]~3_combout ),
	.datad(!\d0_int_bytes_remaining[6]~5_combout ),
	.datae(!\d0_int_bytes_remaining[5]~7_combout ),
	.dataf(!\d0_int_bytes_remaining[4]~8_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\new_burst_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \new_burst_reg~0 .extended_lut = "off";
defparam \new_burst_reg~0 .lut_mask = 64'hAEAAAAAAAAAAAAAA;
defparam \new_burst_reg~0 .shared_arith = "off";

dffeas new_burst_reg(
	.clk(clk_clk),
	.d(\new_burst_reg~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\new_burst_reg~q ),
	.prn(vcc));
defparam new_burst_reg.is_wysiwyg = "true";
defparam new_burst_reg.power_up = "low";

cyclonev_lcell_comb \WideNor0~0 (
	.dataa(!sink0_data[69]),
	.datab(!sink0_data[68]),
	.datac(!WideNor0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideNor0~0 .extended_lut = "off";
defparam \WideNor0~0 .lut_mask = 64'h8A8A8A8A8A8A8A8A;
defparam \WideNor0~0 .shared_arith = "off";

cyclonev_lcell_comb \NON_PIPELINED_INPUTS.load_next_cmd (
	.dataa(!in_ready_hold),
	.datab(!nxt_in_ready1),
	.datac(!nxt_in_ready),
	.datad(!src_valid),
	.datae(!src_valid1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \NON_PIPELINED_INPUTS.load_next_cmd .extended_lut = "off";
defparam \NON_PIPELINED_INPUTS.load_next_cmd .lut_mask = 64'h0015151500151515;
defparam \NON_PIPELINED_INPUTS.load_next_cmd .shared_arith = "off";

dffeas in_bytecount_reg_zero(
	.clk(clk_clk),
	.d(\WideNor0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_bytecount_reg_zero~q ),
	.prn(vcc));
defparam in_bytecount_reg_zero.is_wysiwyg = "true";
defparam in_bytecount_reg_zero.power_up = "low";

cyclonev_lcell_comb \nxt_out_valid~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!\new_burst_reg~q ),
	.datac(!\in_bytecount_reg_zero~q ),
	.datad(!\in_valid~combout ),
	.datae(!cp_ready1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_valid~0 .extended_lut = "off";
defparam \nxt_out_valid~0 .lut_mask = 64'h50FF44FF50FF44FF;
defparam \nxt_out_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!sink0_data[87]),
	.datab(!sink0_data[88]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h8888888888888888;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~0 (
	.dataa(!nxt_out_eop),
	.datab(!\state.ST_UNCOMP_TRANS~q ),
	.datac(!stateST_UNCOMP_WR_SUBBURST),
	.datad(!\WideOr0~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'h002A002A002A002A;
defparam \Selector3~0 .shared_arith = "off";

dffeas \in_size_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[86]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[0]~q ),
	.prn(vcc));
defparam \in_size_reg[0] .is_wysiwyg = "true";
defparam \in_size_reg[0] .power_up = "low";

dffeas \in_size_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[87]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[1]~q ),
	.prn(vcc));
defparam \in_size_reg[1] .is_wysiwyg = "true";
defparam \in_size_reg[1] .power_up = "low";

dffeas \in_size_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[88]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[2]~q ),
	.prn(vcc));
defparam \in_size_reg[2] .is_wysiwyg = "true";
defparam \in_size_reg[2] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[87]),
	.datac(!sink0_data[88]),
	.datad(!\in_size_reg[1]~q ),
	.datae(!\in_size_reg[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~0 .extended_lut = "off";
defparam \ShiftLeft0~0 .lut_mask = 64'h10BA101010BA1010;
defparam \ShiftLeft0~0 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~1 .extended_lut = "off";
defparam \ShiftLeft0~1 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~1 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[3] (
	.clk(clk_clk),
	.d(\ShiftLeft0~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[3]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[3] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[3] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~2 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~2 .extended_lut = "off";
defparam \ShiftLeft0~2 .lut_mask = 64'h00E400E400E400E4;
defparam \ShiftLeft0~2 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[2] (
	.clk(clk_clk),
	.d(\ShiftLeft0~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[2]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[2] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[2] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[87]),
	.datac(!sink0_data[88]),
	.datad(!\in_size_reg[1]~q ),
	.datae(!\in_size_reg[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~3 .extended_lut = "off";
defparam \ShiftLeft0~3 .lut_mask = 64'hEA404040EA404040;
defparam \ShiftLeft0~3 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~4 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~4 .extended_lut = "off";
defparam \ShiftLeft0~4 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~4 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[1] (
	.clk(clk_clk),
	.d(\ShiftLeft0~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[1]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[1] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[1] .power_up = "low";

dffeas \int_byte_cnt_narrow_reg[0] (
	.clk(clk_clk),
	.d(\align_address_to_size|LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[0]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[0] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[0] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[0]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~3 (
	.dataa(!h2f_ARADDR_0),
	.datab(!sink0_data[69]),
	.datac(!sink0_data[68]),
	.datad(!out_data_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~3 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~3 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[0]~3 .shared_arith = "off";

dffeas \in_burstwrap_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[79]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[0]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[0] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[0] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[0]~0 (
	.dataa(!Selector13),
	.datab(!Selector6),
	.datac(!sink0_data[68]),
	.datad(!sink0_data[69]),
	.datae(!\new_burst_reg~q ),
	.dataf(!\d0_int_nxt_addr[0]~4_combout ),
	.datag(!\in_burstwrap_reg[0]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[0]~0 .extended_lut = "on";
defparam \nxt_addr[0]~0 .lut_mask = 64'h00000000F0F0FCA8;
defparam \nxt_addr[0]~0 .shared_arith = "off";

dffeas \int_nxt_addr_reg[0] (
	.clk(clk_clk),
	.d(\nxt_addr[0]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[0] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~4 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\Add0~13_sumout ),
	.datac(!\align_address_to_size|LessThan0~0_combout ),
	.datad(!\d0_int_nxt_addr[0]~3_combout ),
	.datae(!\int_nxt_addr_reg[0]~q ),
	.dataf(!\in_burstwrap_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~4 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~4 .lut_mask = 64'h0005AAAF2227AAAF;
defparam \d0_int_nxt_addr[0]~4 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[0] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[0]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[0] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[1]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[1]~q ),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \in_burstwrap_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[80]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[1]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[1] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[1] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[1]~4 (
	.dataa(!Selector12),
	.datab(!Selector5),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!\new_burst_reg~q ),
	.dataf(!\d0_int_nxt_addr[1]~2_combout ),
	.datag(!\in_burstwrap_reg[1]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[1]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[1]~4 .extended_lut = "on";
defparam \nxt_addr[1]~4 .lut_mask = 64'h00000000F0F0FAC8;
defparam \nxt_addr[1]~4 .shared_arith = "off";

dffeas \int_nxt_addr_reg[1] (
	.clk(clk_clk),
	.d(\nxt_addr[1]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[1] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~7 (
	.dataa(!h2f_ARADDR_1),
	.datab(!sink0_data[69]),
	.datac(!sink0_data[68]),
	.datad(!out_data_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~7 .extended_lut = "off";
defparam \d0_int_nxt_addr[1]~7 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[1]~7 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~2 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\Add0~9_sumout ),
	.datac(!\in_burstwrap_reg[1]~q ),
	.datad(!\int_nxt_addr_reg[1]~q ),
	.datae(!\ShiftLeft0~3_combout ),
	.dataf(!\d0_int_nxt_addr[1]~7_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~2 .extended_lut = "off";
defparam \d0_int_nxt_addr[1]~2 .lut_mask = 64'h02AA02AA02AA57FF;
defparam \d0_int_nxt_addr[1]~2 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[1] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[1]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[1] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_2),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[2]~q ),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[3]~q ),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

dffeas \in_burstwrap_reg[3] (
	.clk(clk_clk),
	.d(sink0_data[82]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[3]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[3] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[3] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[3]~12 (
	.dataa(!Selector10),
	.datab(!Selector3),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!\new_burst_reg~q ),
	.dataf(!\d0_int_nxt_addr[3]~0_combout ),
	.datag(!\in_burstwrap_reg[3]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[3]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[3]~12 .extended_lut = "on";
defparam \nxt_addr[3]~12 .lut_mask = 64'h00000000F0F0FAC8;
defparam \nxt_addr[3]~12 .shared_arith = "off";

dffeas \int_nxt_addr_reg[3] (
	.clk(clk_clk),
	.d(\nxt_addr[3]~12_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[3]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[3] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~5 (
	.dataa(!\Add0~1_sumout ),
	.datab(!\in_burstwrap_reg[3]~q ),
	.datac(!\int_nxt_addr_reg[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~5 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~5 .lut_mask = 64'hE0E0E0E0E0E0E0E0;
defparam \d0_int_nxt_addr[3]~5 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!h2f_ARADDR_3),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!base_address_3),
	.dataf(!\d0_int_nxt_addr[3]~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~0 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~0 .lut_mask = 64'hABABABFF01010155;
defparam \d0_int_nxt_addr[3]~0 .shared_arith = "off";

dffeas \in_burstwrap_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[81]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[2]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[2] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[2] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[2]~8 (
	.dataa(!Selector11),
	.datab(!Selector4),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!\new_burst_reg~q ),
	.dataf(!\d0_int_nxt_addr[2]~1_combout ),
	.datag(!\in_burstwrap_reg[2]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[2]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[2]~8 .extended_lut = "on";
defparam \nxt_addr[2]~8 .lut_mask = 64'h00000000F0F0FAC8;
defparam \nxt_addr[2]~8 .shared_arith = "off";

dffeas \int_nxt_addr_reg[2] (
	.clk(clk_clk),
	.d(\nxt_addr[2]~8_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[2]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~6 (
	.dataa(!\Add0~5_sumout ),
	.datab(!\in_burstwrap_reg[2]~q ),
	.datac(!\int_nxt_addr_reg[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~6 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~6 .lut_mask = 64'hE0E0E0E0E0E0E0E0;
defparam \d0_int_nxt_addr[2]~6 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!h2f_ARADDR_2),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!base_address_2),
	.dataf(!\d0_int_nxt_addr[2]~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~1 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~1 .lut_mask = 64'hABABABFF01010155;
defparam \d0_int_nxt_addr[2]~1 .shared_arith = "off";

dffeas in_eop_reg(
	.clk(clk_clk),
	.d(sink0_endofpacket),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_eop_reg~q ),
	.prn(vcc));
defparam in_eop_reg.is_wysiwyg = "true";
defparam in_eop_reg.power_up = "low";

endmodule

module spw_babasu_altera_merlin_address_alignment_3 (
	new_burst_reg,
	src_data_86,
	in_size_reg_0,
	ShiftLeft0,
	LessThan0)/* synthesis synthesis_greybox=0 */;
input 	new_burst_reg;
input 	src_data_86;
input 	in_size_reg_0;
input 	ShiftLeft0;
output 	LessThan0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!new_burst_reg),
	.datab(!src_data_86),
	.datac(!in_size_reg_0),
	.datad(!ShiftLeft0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan0),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h00E400E400E400E4;
defparam \LessThan0~0 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_burst_adapter_3 (
	h2f_ARADDR_0,
	h2f_ARADDR_1,
	h2f_ARADDR_2,
	h2f_ARADDR_3,
	h2f_ARBURST_0,
	h2f_ARBURST_1,
	h2f_ARID_0,
	h2f_ARID_1,
	h2f_ARID_2,
	h2f_ARID_3,
	h2f_ARID_4,
	h2f_ARID_5,
	h2f_ARID_6,
	h2f_ARID_7,
	h2f_ARID_8,
	h2f_ARID_9,
	h2f_ARID_10,
	h2f_ARID_11,
	h2f_ARLEN_0,
	Add5,
	Add51,
	saved_grant_1,
	stateST_COMP_TRANS,
	mem_used_1,
	in_data_reg_69,
	in_narrow_reg,
	cp_ready,
	cp_ready1,
	nxt_out_eop,
	in_ready_hold,
	out_valid_reg,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready,
	altera_reset_synchronizer_int_chain_out,
	nxt_in_ready1,
	src_valid,
	Decoder1,
	out_byte_cnt_reg_2,
	Add2,
	Add21,
	Add22,
	Add23,
	cp_ready2,
	out_uncomp_byte_cnt_reg_6,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	Selector10,
	Selector101,
	Selector11,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	Selector12,
	src_payload,
	src_payload1,
	src_payload2,
	Selector13,
	nxt_out_burstwrap_1,
	nxt_addr_2,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARADDR_0;
input 	h2f_ARADDR_1;
input 	h2f_ARADDR_2;
input 	h2f_ARADDR_3;
input 	h2f_ARBURST_0;
input 	h2f_ARBURST_1;
input 	h2f_ARID_0;
input 	h2f_ARID_1;
input 	h2f_ARID_2;
input 	h2f_ARID_3;
input 	h2f_ARID_4;
input 	h2f_ARID_5;
input 	h2f_ARID_6;
input 	h2f_ARID_7;
input 	h2f_ARID_8;
input 	h2f_ARID_9;
input 	h2f_ARID_10;
input 	h2f_ARID_11;
input 	h2f_ARLEN_0;
input 	Add5;
input 	Add51;
input 	saved_grant_1;
output 	stateST_COMP_TRANS;
input 	mem_used_1;
output 	in_data_reg_69;
output 	in_narrow_reg;
input 	cp_ready;
input 	cp_ready1;
output 	nxt_out_eop;
input 	in_ready_hold;
output 	out_valid_reg;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready;
input 	altera_reset_synchronizer_int_chain_out;
output 	nxt_in_ready1;
input 	src_valid;
input 	Decoder1;
output 	out_byte_cnt_reg_2;
input 	Add2;
input 	Add21;
input 	Add22;
input 	Add23;
input 	cp_ready2;
output 	out_uncomp_byte_cnt_reg_6;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	in_data_reg_105;
output 	in_data_reg_106;
output 	in_data_reg_107;
output 	in_data_reg_108;
output 	in_data_reg_109;
output 	in_data_reg_110;
output 	in_data_reg_111;
output 	in_data_reg_112;
output 	in_data_reg_113;
output 	in_data_reg_114;
output 	in_data_reg_115;
output 	in_data_reg_116;
input 	Selector10;
input 	Selector101;
input 	Selector11;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
input 	Selector12;
input 	src_payload;
input 	src_payload1;
input 	src_payload2;
input 	Selector13;
input 	nxt_out_burstwrap_1;
input 	nxt_addr_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



spw_babasu_altera_merlin_burst_adapter_13_1_3 \altera_merlin_burst_adapter_13_1.burst_adapter (
	.h2f_ARADDR_0(h2f_ARADDR_0),
	.h2f_ARADDR_1(h2f_ARADDR_1),
	.h2f_ARADDR_2(h2f_ARADDR_2),
	.h2f_ARADDR_3(h2f_ARADDR_3),
	.h2f_ARBURST_0(h2f_ARBURST_0),
	.h2f_ARBURST_1(h2f_ARBURST_1),
	.sink0_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,h2f_ARID_11,h2f_ARID_10,h2f_ARID_9,h2f_ARID_8,h2f_ARID_7,h2f_ARID_6,h2f_ARID_5,h2f_ARID_4,h2f_ARID_3,h2f_ARID_2,h2f_ARID_1,h2f_ARID_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_payload1,src_payload2,src_payload,gnd,gnd,gnd,
Selector101,Selector11,Selector12,Selector13,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,saved_grant_1,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.h2f_ARLEN_0(h2f_ARLEN_0),
	.Add5(Add5),
	.Add51(Add51),
	.stateST_COMP_TRANS(stateST_COMP_TRANS),
	.mem_used_1(mem_used_1),
	.in_data_reg_69(in_data_reg_69),
	.in_narrow_reg1(in_narrow_reg),
	.cp_ready(cp_ready),
	.cp_ready1(cp_ready1),
	.nxt_out_eop(nxt_out_eop),
	.in_ready_hold(in_ready_hold),
	.out_valid_reg1(out_valid_reg),
	.stateST_UNCOMP_WR_SUBBURST(stateST_UNCOMP_WR_SUBBURST),
	.nxt_in_ready(nxt_in_ready),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.nxt_in_ready1(nxt_in_ready1),
	.src_valid(src_valid),
	.Decoder1(Decoder1),
	.out_byte_cnt_reg_2(out_byte_cnt_reg_2),
	.Add2(Add2),
	.Add21(Add21),
	.Add22(Add22),
	.Add23(Add23),
	.cp_ready2(cp_ready2),
	.out_uncomp_byte_cnt_reg_6(out_uncomp_byte_cnt_reg_6),
	.out_uncomp_byte_cnt_reg_5(out_uncomp_byte_cnt_reg_5),
	.out_uncomp_byte_cnt_reg_4(out_uncomp_byte_cnt_reg_4),
	.out_uncomp_byte_cnt_reg_3(out_uncomp_byte_cnt_reg_3),
	.out_uncomp_byte_cnt_reg_2(out_uncomp_byte_cnt_reg_2),
	.in_data_reg_105(in_data_reg_105),
	.in_data_reg_106(in_data_reg_106),
	.in_data_reg_107(in_data_reg_107),
	.in_data_reg_108(in_data_reg_108),
	.in_data_reg_109(in_data_reg_109),
	.in_data_reg_110(in_data_reg_110),
	.in_data_reg_111(in_data_reg_111),
	.in_data_reg_112(in_data_reg_112),
	.in_data_reg_113(in_data_reg_113),
	.in_data_reg_114(in_data_reg_114),
	.in_data_reg_115(in_data_reg_115),
	.in_data_reg_116(in_data_reg_116),
	.Selector10(Selector10),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_3),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_2),
	.nxt_out_burstwrap_1(nxt_out_burstwrap_1),
	.nxt_addr_2(nxt_addr_2),
	.clk_clk(clk_clk));

endmodule

module spw_babasu_altera_merlin_burst_adapter_13_1_3 (
	h2f_ARADDR_0,
	h2f_ARADDR_1,
	h2f_ARADDR_2,
	h2f_ARADDR_3,
	h2f_ARBURST_0,
	h2f_ARBURST_1,
	sink0_data,
	h2f_ARLEN_0,
	Add5,
	Add51,
	stateST_COMP_TRANS,
	mem_used_1,
	in_data_reg_69,
	in_narrow_reg1,
	cp_ready,
	cp_ready1,
	nxt_out_eop,
	in_ready_hold,
	out_valid_reg1,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready,
	altera_reset_synchronizer_int_chain_out,
	nxt_in_ready1,
	src_valid,
	Decoder1,
	out_byte_cnt_reg_2,
	Add2,
	Add21,
	Add22,
	Add23,
	cp_ready2,
	out_uncomp_byte_cnt_reg_6,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	Selector10,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	nxt_out_burstwrap_1,
	nxt_addr_2,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARADDR_0;
input 	h2f_ARADDR_1;
input 	h2f_ARADDR_2;
input 	h2f_ARADDR_3;
input 	h2f_ARBURST_0;
input 	h2f_ARBURST_1;
input 	[128:0] sink0_data;
input 	h2f_ARLEN_0;
input 	Add5;
input 	Add51;
output 	stateST_COMP_TRANS;
input 	mem_used_1;
output 	in_data_reg_69;
output 	in_narrow_reg1;
input 	cp_ready;
input 	cp_ready1;
output 	nxt_out_eop;
input 	in_ready_hold;
output 	out_valid_reg1;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready;
input 	altera_reset_synchronizer_int_chain_out;
output 	nxt_in_ready1;
input 	src_valid;
input 	Decoder1;
output 	out_byte_cnt_reg_2;
input 	Add2;
input 	Add21;
input 	Add22;
input 	Add23;
input 	cp_ready2;
output 	out_uncomp_byte_cnt_reg_6;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	in_data_reg_105;
output 	in_data_reg_106;
output 	in_data_reg_107;
output 	in_data_reg_108;
output 	in_data_reg_109;
output 	in_data_reg_110;
output 	in_data_reg_111;
output 	in_data_reg_112;
output 	in_data_reg_113;
output 	in_data_reg_114;
output 	in_data_reg_115;
output 	in_data_reg_116;
input 	Selector10;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
input 	nxt_out_burstwrap_1;
input 	nxt_addr_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \align_address_to_size|LessThan0~0_combout ;
wire \align_address_to_size|LessThan0~1_combout ;
wire \nxt_uncomp_subburst_byte_cnt~0_combout ;
wire \Add4~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt[6]~1_combout ;
wire \nxt_uncomp_subburst_byte_cnt[5]~2_combout ;
wire \nxt_uncomp_subburst_byte_cnt[4]~3_combout ;
wire \nxt_uncomp_subburst_byte_cnt[3]~4_combout ;
wire \nxt_uncomp_subburst_byte_cnt[2]~5_combout ;
wire \WideNor1~combout ;
wire \Selector2~1_combout ;
wire \load_next_out_cmd~combout ;
wire \state.ST_UNCOMP_TRANS~q ;
wire \Selector2~0_combout ;
wire \Selector0~0_combout ;
wire \state.ST_IDLE~q ;
wire \Selector1~0_combout ;
wire \Selector1~1_combout ;
wire \NON_PIPELINED_INPUTS.load_next_cmd~0_combout ;
wire \int_bytes_remaining_reg[2]~q ;
wire \d0_int_bytes_remaining[2]~0_combout ;
wire \int_bytes_remaining_reg[3]~q ;
wire \d0_int_bytes_remaining[3]~1_combout ;
wire \int_bytes_remaining_reg[4]~q ;
wire \Add1~0_combout ;
wire \d0_int_bytes_remaining[4]~2_combout ;
wire \int_bytes_remaining_reg[5]~q ;
wire \Add1~1_combout ;
wire \d0_int_bytes_remaining[5]~3_combout ;
wire \int_bytes_remaining_reg[6]~q ;
wire \d0_int_bytes_remaining[6]~4_combout ;
wire \new_burst_reg~0_combout ;
wire \new_burst_reg~q ;
wire \in_bytecount_reg_zero~0_combout ;
wire \in_bytecount_reg_zero~q ;
wire \nxt_out_valid~0_combout ;
wire \nxt_out_valid~1_combout ;
wire \Selector3~0_combout ;
wire \in_burstwrap_reg[3]~q ;
wire \nxt_addr[3]~0_combout ;
wire \nxt_addr[3]~combout ;
wire \int_nxt_addr_reg[3]~q ;
wire \in_size_reg[0]~q ;
wire \in_size_reg[2]~q ;
wire \in_size_reg[1]~q ;
wire \ShiftLeft0~0_combout ;
wire \ShiftLeft0~1_combout ;
wire \int_byte_cnt_narrow_reg[3]~q ;
wire \ShiftLeft0~2_combout ;
wire \int_byte_cnt_narrow_reg[2]~q ;
wire \in_burstwrap_reg[1]~q ;
wire \nxt_addr[1]~combout ;
wire \int_nxt_addr_reg[1]~q ;
wire \ShiftLeft0~3_combout ;
wire \int_byte_cnt_narrow_reg[1]~q ;
wire \int_byte_cnt_narrow_reg[0]~q ;
wire \Add0~13_sumout ;
wire \in_burstwrap_reg[0]~q ;
wire \nxt_addr[0]~combout ;
wire \int_nxt_addr_reg[0]~q ;
wire \d0_int_nxt_addr[0]~2_combout ;
wire \d0_int_nxt_addr[0]~3_combout ;
wire \int_nxt_addr_reg_dly[0]~q ;
wire \Add0~14 ;
wire \Add0~9_sumout ;
wire \d0_int_nxt_addr[1]~4_combout ;
wire \int_nxt_addr_reg_dly[1]~q ;
wire \Add0~10 ;
wire \Add0~6 ;
wire \Add0~1_sumout ;
wire \d0_int_nxt_addr[3]~0_combout ;
wire \in_burstwrap_reg[2]~q ;
wire \nxt_addr[2]~1_combout ;
wire \nxt_addr[2]~combout ;
wire \int_nxt_addr_reg[2]~q ;
wire \Add0~5_sumout ;
wire \d0_int_nxt_addr[2]~1_combout ;


spw_babasu_altera_merlin_address_alignment_4 align_address_to_size(
	.new_burst_reg(\new_burst_reg~q ),
	.src_payload(sink0_data[86]),
	.in_size_reg_0(\in_size_reg[0]~q ),
	.src_payload1(sink0_data[88]),
	.in_size_reg_2(\in_size_reg[2]~q ),
	.src_payload2(sink0_data[87]),
	.in_size_reg_1(\in_size_reg[1]~q ),
	.LessThan0(\align_address_to_size|LessThan0~0_combout ),
	.LessThan01(\align_address_to_size|LessThan0~1_combout ));

dffeas \state.ST_COMP_TRANS (
	.clk(clk_clk),
	.d(\Selector1~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_COMP_TRANS),
	.prn(vcc));
defparam \state.ST_COMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_COMP_TRANS .power_up = "low";

dffeas \in_data_reg[69] (
	.clk(clk_clk),
	.d(sink0_data[69]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_69),
	.prn(vcc));
defparam \in_data_reg[69] .is_wysiwyg = "true";
defparam \in_data_reg[69] .power_up = "low";

dffeas in_narrow_reg(
	.clk(clk_clk),
	.d(Decoder1),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_narrow_reg1),
	.prn(vcc));
defparam in_narrow_reg.is_wysiwyg = "true";
defparam in_narrow_reg.power_up = "low";

cyclonev_lcell_comb \nxt_out_eop~0 (
	.dataa(!in_data_reg_69),
	.datab(!stateST_COMP_TRANS),
	.datac(!\new_burst_reg~q ),
	.datad(!mem_used_1),
	.datae(!cp_ready),
	.dataf(!\in_bytecount_reg_zero~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_out_eop),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_eop~0 .extended_lut = "off";
defparam \nxt_out_eop~0 .lut_mask = 64'h4444474477774777;
defparam \nxt_out_eop~0 .shared_arith = "off";

dffeas out_valid_reg(
	.clk(clk_clk),
	.d(\nxt_out_valid~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_valid_reg1),
	.prn(vcc));
defparam out_valid_reg.is_wysiwyg = "true";
defparam out_valid_reg.power_up = "low";

dffeas \state.ST_UNCOMP_WR_SUBBURST (
	.clk(clk_clk),
	.d(\Selector3~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_UNCOMP_WR_SUBBURST),
	.prn(vcc));
defparam \state.ST_UNCOMP_WR_SUBBURST .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_WR_SUBBURST .power_up = "low";

cyclonev_lcell_comb \nxt_in_ready~0 (
	.dataa(!in_ready_hold),
	.datab(!stateST_COMP_TRANS),
	.datac(!mem_used_1),
	.datad(!cp_ready),
	.datae(!out_valid_reg1),
	.dataf(!\Selector2~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~0 .extended_lut = "off";
defparam \nxt_in_ready~0 .lut_mask = 64'h0000FF3F8888BBBB;
defparam \nxt_in_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_in_ready~1 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!cp_ready1),
	.datac(!nxt_out_eop),
	.datad(!nxt_in_ready),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~1 .extended_lut = "off";
defparam \nxt_in_ready~1 .lut_mask = 64'h00FE00FE00FE00FE;
defparam \nxt_in_ready~1 .shared_arith = "off";

dffeas \out_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[6] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[6]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_6),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[6] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[6] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[5] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[5]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_5),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[5] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[5] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[4] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[4]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_4),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[4] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[4] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[3] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[3]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_3),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[3] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[3] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[2]~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[2] .power_up = "low";

dffeas \in_data_reg[105] (
	.clk(clk_clk),
	.d(sink0_data[105]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_105),
	.prn(vcc));
defparam \in_data_reg[105] .is_wysiwyg = "true";
defparam \in_data_reg[105] .power_up = "low";

dffeas \in_data_reg[106] (
	.clk(clk_clk),
	.d(sink0_data[106]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_106),
	.prn(vcc));
defparam \in_data_reg[106] .is_wysiwyg = "true";
defparam \in_data_reg[106] .power_up = "low";

dffeas \in_data_reg[107] (
	.clk(clk_clk),
	.d(sink0_data[107]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_107),
	.prn(vcc));
defparam \in_data_reg[107] .is_wysiwyg = "true";
defparam \in_data_reg[107] .power_up = "low";

dffeas \in_data_reg[108] (
	.clk(clk_clk),
	.d(sink0_data[108]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_108),
	.prn(vcc));
defparam \in_data_reg[108] .is_wysiwyg = "true";
defparam \in_data_reg[108] .power_up = "low";

dffeas \in_data_reg[109] (
	.clk(clk_clk),
	.d(sink0_data[109]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_109),
	.prn(vcc));
defparam \in_data_reg[109] .is_wysiwyg = "true";
defparam \in_data_reg[109] .power_up = "low";

dffeas \in_data_reg[110] (
	.clk(clk_clk),
	.d(sink0_data[110]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_110),
	.prn(vcc));
defparam \in_data_reg[110] .is_wysiwyg = "true";
defparam \in_data_reg[110] .power_up = "low";

dffeas \in_data_reg[111] (
	.clk(clk_clk),
	.d(sink0_data[111]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_111),
	.prn(vcc));
defparam \in_data_reg[111] .is_wysiwyg = "true";
defparam \in_data_reg[111] .power_up = "low";

dffeas \in_data_reg[112] (
	.clk(clk_clk),
	.d(sink0_data[112]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_112),
	.prn(vcc));
defparam \in_data_reg[112] .is_wysiwyg = "true";
defparam \in_data_reg[112] .power_up = "low";

dffeas \in_data_reg[113] (
	.clk(clk_clk),
	.d(sink0_data[113]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_113),
	.prn(vcc));
defparam \in_data_reg[113] .is_wysiwyg = "true";
defparam \in_data_reg[113] .power_up = "low";

dffeas \in_data_reg[114] (
	.clk(clk_clk),
	.d(sink0_data[114]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_114),
	.prn(vcc));
defparam \in_data_reg[114] .is_wysiwyg = "true";
defparam \in_data_reg[114] .power_up = "low";

dffeas \in_data_reg[115] (
	.clk(clk_clk),
	.d(sink0_data[115]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_115),
	.prn(vcc));
defparam \in_data_reg[115] .is_wysiwyg = "true";
defparam \in_data_reg[115] .power_up = "low";

dffeas \in_data_reg[116] (
	.clk(clk_clk),
	.d(sink0_data[116]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_116),
	.prn(vcc));
defparam \in_data_reg[116] .is_wysiwyg = "true";
defparam \in_data_reg[116] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[3] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[3]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_3),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[3] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[2] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[2]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_2),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[2] .power_up = "low";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt~0 (
	.dataa(!cp_ready1),
	.datab(!out_valid_reg1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt~0 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt~0 .lut_mask = 64'h1111111111111111;
defparam \nxt_uncomp_subburst_byte_cnt~0 .shared_arith = "off";

cyclonev_lcell_comb \Add4~0 (
	.dataa(!out_uncomp_byte_cnt_reg_4),
	.datab(!out_uncomp_byte_cnt_reg_3),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add4~0 .extended_lut = "off";
defparam \Add4~0 .lut_mask = 64'h0800080008000800;
defparam \Add4~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[6]~1 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_6),
	.datad(!out_uncomp_byte_cnt_reg_5),
	.datae(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.dataf(!\Add4~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[6]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[6]~1 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[6]~1 .lut_mask = 64'h0F0F4E4EA50FE44E;
defparam \nxt_uncomp_subburst_byte_cnt[6]~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[5]~2 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!\Add4~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[5]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[5]~2 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[5]~2 .lut_mask = 64'h0F4EA5E40F4EA5E4;
defparam \nxt_uncomp_subburst_byte_cnt[5]~2 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[4]~3 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!out_uncomp_byte_cnt_reg_3),
	.datae(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.dataf(!out_uncomp_byte_cnt_reg_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[4]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[4]~3 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[4]~3 .lut_mask = 64'h0F0FE44E0F0F4E4E;
defparam \nxt_uncomp_subburst_byte_cnt[4]~3 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[3]~4 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!out_uncomp_byte_cnt_reg_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[3]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[3]~4 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[3]~4 .lut_mask = 64'h0FE40F4E0FE40F4E;
defparam \nxt_uncomp_subburst_byte_cnt[3]~4 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[2]~5 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[2]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[2]~5 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[2]~5 .lut_mask = 64'h0EF40EF40EF40EF4;
defparam \nxt_uncomp_subburst_byte_cnt[2]~5 .shared_arith = "off";

cyclonev_lcell_comb WideNor1(
	.dataa(!\nxt_uncomp_subburst_byte_cnt[6]~1_combout ),
	.datab(!\nxt_uncomp_subburst_byte_cnt[5]~2_combout ),
	.datac(!\nxt_uncomp_subburst_byte_cnt[4]~3_combout ),
	.datad(!\nxt_uncomp_subburst_byte_cnt[3]~4_combout ),
	.datae(!\nxt_uncomp_subburst_byte_cnt[2]~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideNor1.extended_lut = "off";
defparam WideNor1.lut_mask = 64'h8000000080000000;
defparam WideNor1.shared_arith = "off";

cyclonev_lcell_comb \Selector2~1 (
	.dataa(!nxt_out_eop),
	.datab(!\Selector2~0_combout ),
	.datac(!\WideNor1~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~1 .extended_lut = "off";
defparam \Selector2~1 .lut_mask = 64'h0808080808080808;
defparam \Selector2~1 .shared_arith = "off";

cyclonev_lcell_comb load_next_out_cmd(
	.dataa(!mem_used_1),
	.datab(!cp_ready),
	.datac(!out_valid_reg1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\load_next_out_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam load_next_out_cmd.extended_lut = "off";
defparam load_next_out_cmd.lut_mask = 64'hF2F2F2F2F2F2F2F2;
defparam load_next_out_cmd.shared_arith = "off";

dffeas \state.ST_UNCOMP_TRANS (
	.clk(clk_clk),
	.d(\Selector2~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_UNCOMP_TRANS~q ),
	.prn(vcc));
defparam \state.ST_UNCOMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_TRANS .power_up = "low";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'h8888888888888888;
defparam \Selector2~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!in_ready_hold),
	.datab(!nxt_out_eop),
	.datac(!src_valid),
	.datad(!\state.ST_IDLE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'h05CD05CD05CD05CD;
defparam \Selector0~0 .shared_arith = "off";

dffeas \state.ST_IDLE (
	.clk(clk_clk),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_IDLE~q ),
	.prn(vcc));
defparam \state.ST_IDLE .is_wysiwyg = "true";
defparam \state.ST_IDLE .power_up = "low";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!sink0_data[69]),
	.datab(!nxt_out_eop),
	.datac(!\Selector2~0_combout ),
	.datad(!\state.ST_IDLE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'h5510551055105510;
defparam \Selector1~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~1 (
	.dataa(!in_ready_hold),
	.datab(!stateST_COMP_TRANS),
	.datac(!nxt_out_eop),
	.datad(!src_valid),
	.datae(!\Selector1~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~1 .extended_lut = "off";
defparam \Selector1~1 .lut_mask = 64'h3031307530313075;
defparam \Selector1~1 .shared_arith = "off";

cyclonev_lcell_comb \NON_PIPELINED_INPUTS.load_next_cmd~0 (
	.dataa(!in_ready_hold),
	.datab(!nxt_in_ready1),
	.datac(!src_valid),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \NON_PIPELINED_INPUTS.load_next_cmd~0 .extended_lut = "off";
defparam \NON_PIPELINED_INPUTS.load_next_cmd~0 .lut_mask = 64'h0404040404040404;
defparam \NON_PIPELINED_INPUTS.load_next_cmd~0 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[2] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[2]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[2]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[2] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[2]~0 (
	.dataa(!h2f_ARLEN_0),
	.datab(!sink0_data[69]),
	.datac(!\new_burst_reg~q ),
	.datad(!out_byte_cnt_reg_2),
	.datae(!\int_bytes_remaining_reg[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[2]~0 .extended_lut = "off";
defparam \d0_int_bytes_remaining[2]~0 .lut_mask = 64'h02F2F20202F2F202;
defparam \d0_int_bytes_remaining[2]~0 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[3] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[3]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[3]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[3] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[3] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[3]~1 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!Add2),
	.datad(!out_byte_cnt_reg_2),
	.datae(!\int_bytes_remaining_reg[2]~q ),
	.dataf(!\int_bytes_remaining_reg[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[3]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[3]~1 .extended_lut = "off";
defparam \d0_int_bytes_remaining[3]~1 .lut_mask = 64'h01CD0101CD01CDCD;
defparam \d0_int_bytes_remaining[3]~1 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[4] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[4]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[4]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[4] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[4] .power_up = "low";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!out_byte_cnt_reg_2),
	.datab(!\int_bytes_remaining_reg[2]~q ),
	.datac(!\int_bytes_remaining_reg[3]~q ),
	.datad(!\int_bytes_remaining_reg[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'hBF40BF40BF40BF40;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[4]~2 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!Add21),
	.datad(!\Add1~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[4]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[4]~2 .extended_lut = "off";
defparam \d0_int_bytes_remaining[4]~2 .lut_mask = 64'hCD01CD01CD01CD01;
defparam \d0_int_bytes_remaining[4]~2 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[5] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[5]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[5]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[5] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[5] .power_up = "low";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!out_byte_cnt_reg_2),
	.datab(!\int_bytes_remaining_reg[2]~q ),
	.datac(!\int_bytes_remaining_reg[3]~q ),
	.datad(!\int_bytes_remaining_reg[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h4000400040004000;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[5]~3 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!Add22),
	.datad(!\int_bytes_remaining_reg[5]~q ),
	.datae(!\Add1~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[5]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[5]~3 .extended_lut = "off";
defparam \d0_int_bytes_remaining[5]~3 .lut_mask = 64'h01CDCD0101CDCD01;
defparam \d0_int_bytes_remaining[5]~3 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[6] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[6]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[6]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[6] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[6] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[6]~4 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!Add23),
	.datad(!\int_bytes_remaining_reg[5]~q ),
	.datae(!\Add1~1_combout ),
	.dataf(!\int_bytes_remaining_reg[6]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[6]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[6]~4 .extended_lut = "off";
defparam \d0_int_bytes_remaining[6]~4 .lut_mask = 64'h0101CD01CDCD01CD;
defparam \d0_int_bytes_remaining[6]~4 .shared_arith = "off";

cyclonev_lcell_comb \new_burst_reg~0 (
	.dataa(!\Selector1~1_combout ),
	.datab(!\d0_int_bytes_remaining[2]~0_combout ),
	.datac(!\d0_int_bytes_remaining[3]~1_combout ),
	.datad(!\d0_int_bytes_remaining[4]~2_combout ),
	.datae(!\d0_int_bytes_remaining[5]~3_combout ),
	.dataf(!\d0_int_bytes_remaining[6]~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\new_burst_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \new_burst_reg~0 .extended_lut = "off";
defparam \new_burst_reg~0 .lut_mask = 64'hBAAAAAAAAAAAAAAA;
defparam \new_burst_reg~0 .shared_arith = "off";

dffeas new_burst_reg(
	.clk(clk_clk),
	.d(\new_burst_reg~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\new_burst_reg~q ),
	.prn(vcc));
defparam new_burst_reg.is_wysiwyg = "true";
defparam new_burst_reg.power_up = "low";

cyclonev_lcell_comb \in_bytecount_reg_zero~0 (
	.dataa(!sink0_data[69]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\in_bytecount_reg_zero~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \in_bytecount_reg_zero~0 .extended_lut = "off";
defparam \in_bytecount_reg_zero~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \in_bytecount_reg_zero~0 .shared_arith = "off";

dffeas in_bytecount_reg_zero(
	.clk(clk_clk),
	.d(\in_bytecount_reg_zero~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_bytecount_reg_zero~q ),
	.prn(vcc));
defparam in_bytecount_reg_zero.is_wysiwyg = "true";
defparam in_bytecount_reg_zero.power_up = "low";

cyclonev_lcell_comb \nxt_out_valid~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!mem_used_1),
	.datac(!\in_bytecount_reg_zero~q ),
	.datad(!cp_ready2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_valid~0 .extended_lut = "off";
defparam \nxt_out_valid~0 .lut_mask = 64'hF0B8F0B8F0B8F0B8;
defparam \nxt_out_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_out_valid~1 (
	.dataa(!in_ready_hold),
	.datab(!stateST_COMP_TRANS),
	.datac(!src_valid),
	.datad(!\nxt_out_valid~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_valid~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_valid~1 .extended_lut = "off";
defparam \nxt_out_valid~1 .lut_mask = 64'h0537053705370537;
defparam \nxt_out_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~0 (
	.dataa(!nxt_out_eop),
	.datab(!\Selector2~0_combout ),
	.datac(!\WideNor1~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'h8080808080808080;
defparam \Selector3~0 .shared_arith = "off";

dffeas \in_burstwrap_reg[3] (
	.clk(clk_clk),
	.d(sink0_data[82]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_burstwrap_reg[3]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[3] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[3] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[3]~0 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!\in_burstwrap_reg[3]~q ),
	.datad(!\d0_int_nxt_addr[3]~0_combout ),
	.datae(!h2f_ARBURST_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[3]~0 .extended_lut = "off";
defparam \nxt_addr[3]~0 .lut_mask = 64'h00F300E200F300E2;
defparam \nxt_addr[3]~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_addr[3] (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!h2f_ARBURST_1),
	.datad(!Add5),
	.datae(!Selector10),
	.dataf(!\nxt_addr[3]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[3] .extended_lut = "off";
defparam \nxt_addr[3] .lut_mask = 64'h00000000FEEEFFEF;
defparam \nxt_addr[3] .shared_arith = "off";

dffeas \int_nxt_addr_reg[3] (
	.clk(clk_clk),
	.d(\nxt_addr[3]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[3]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[3] .power_up = "low";

dffeas \in_size_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[86]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_size_reg[0]~q ),
	.prn(vcc));
defparam \in_size_reg[0] .is_wysiwyg = "true";
defparam \in_size_reg[0] .power_up = "low";

dffeas \in_size_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[88]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_size_reg[2]~q ),
	.prn(vcc));
defparam \in_size_reg[2] .is_wysiwyg = "true";
defparam \in_size_reg[2] .power_up = "low";

dffeas \in_size_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[87]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_size_reg[1]~q ),
	.prn(vcc));
defparam \in_size_reg[1] .is_wysiwyg = "true";
defparam \in_size_reg[1] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[88]),
	.datac(!\in_size_reg[2]~q ),
	.datad(!sink0_data[87]),
	.datae(!\in_size_reg[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~0 .extended_lut = "off";
defparam \ShiftLeft0~0 .lut_mask = 64'h0044A0E40044A0E4;
defparam \ShiftLeft0~0 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~1 .extended_lut = "off";
defparam \ShiftLeft0~1 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~1 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[3] (
	.clk(clk_clk),
	.d(\ShiftLeft0~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[3]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[3] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[3] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~2 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~2 .extended_lut = "off";
defparam \ShiftLeft0~2 .lut_mask = 64'h00E400E400E400E4;
defparam \ShiftLeft0~2 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[2] (
	.clk(clk_clk),
	.d(\ShiftLeft0~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[2]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[2] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[2] .power_up = "low";

dffeas \in_burstwrap_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[80]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_burstwrap_reg[1]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[1] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[1] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[1] (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!\in_burstwrap_reg[1]~q ),
	.datad(!\d0_int_nxt_addr[1]~4_combout ),
	.datae(!nxt_out_burstwrap_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[1] .extended_lut = "off";
defparam \nxt_addr[1] .lut_mask = 64'h00E200F300E200F3;
defparam \nxt_addr[1] .shared_arith = "off";

dffeas \int_nxt_addr_reg[1] (
	.clk(clk_clk),
	.d(\nxt_addr[1]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[1] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\align_address_to_size|LessThan0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~3 .extended_lut = "off";
defparam \ShiftLeft0~3 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~3 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[1] (
	.clk(clk_clk),
	.d(\ShiftLeft0~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[1]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[1] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[1] .power_up = "low";

dffeas \int_byte_cnt_narrow_reg[0] (
	.clk(clk_clk),
	.d(\align_address_to_size|LessThan0~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[0]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[0] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[0] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[0]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \in_burstwrap_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[79]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_burstwrap_reg[0]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[0] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[0] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[0] (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!sink0_data[79]),
	.datad(!\in_burstwrap_reg[0]~q ),
	.datae(!\d0_int_nxt_addr[0]~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[0] .extended_lut = "off";
defparam \nxt_addr[0] .lut_mask = 64'h0000FE320000FE32;
defparam \nxt_addr[0] .shared_arith = "off";

dffeas \int_nxt_addr_reg[0] (
	.clk(clk_clk),
	.d(\nxt_addr[0]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[0] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~2 (
	.dataa(!\Add0~13_sumout ),
	.datab(!\int_nxt_addr_reg[0]~q ),
	.datac(!\in_burstwrap_reg[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~2 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~2 .lut_mask = 64'hC8C8C8C8C8C8C8C8;
defparam \d0_int_nxt_addr[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~3 (
	.dataa(!h2f_ARADDR_0),
	.datab(!sink0_data[69]),
	.datac(!\new_burst_reg~q ),
	.datad(!\align_address_to_size|LessThan0~1_combout ),
	.datae(!\d0_int_nxt_addr[0]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~3 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~3 .lut_mask = 64'hF0F10001F0F10001;
defparam \d0_int_nxt_addr[0]~3 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[0] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[0]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[0] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[1]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[1]~q ),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~4 (
	.dataa(!\int_nxt_addr_reg[1]~q ),
	.datab(!\Add0~9_sumout ),
	.datac(!sink0_data[69]),
	.datad(!Decoder1),
	.datae(!\new_burst_reg~q ),
	.dataf(!h2f_ARADDR_1),
	.datag(!\in_burstwrap_reg[1]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~4 .extended_lut = "on";
defparam \d0_int_nxt_addr[1]~4 .lut_mask = 64'h575700005757000F;
defparam \d0_int_nxt_addr[1]~4 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[1] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[1]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[1] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_2),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[2]~q ),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[3]~q ),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~0 (
	.dataa(!h2f_ARADDR_3),
	.datab(!sink0_data[69]),
	.datac(!\new_burst_reg~q ),
	.datad(!\int_nxt_addr_reg[3]~q ),
	.datae(!\in_burstwrap_reg[3]~q ),
	.dataf(!\Add0~1_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~0 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~0 .lut_mask = 64'h01F101F101F1F1F1;
defparam \d0_int_nxt_addr[3]~0 .shared_arith = "off";

dffeas \in_burstwrap_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[81]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_burstwrap_reg[2]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[2] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[2] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[2]~1 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!\in_burstwrap_reg[2]~q ),
	.datad(!\d0_int_nxt_addr[2]~1_combout ),
	.datae(!h2f_ARBURST_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[2]~1 .extended_lut = "off";
defparam \nxt_addr[2]~1 .lut_mask = 64'h00F300E200F300E2;
defparam \nxt_addr[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_addr[2] (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!h2f_ARBURST_1),
	.datad(!Add51),
	.datae(!\nxt_addr[2]~1_combout ),
	.dataf(!nxt_addr_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[2] .extended_lut = "off";
defparam \nxt_addr[2] .lut_mask = 64'h0000FEEE0000FFEF;
defparam \nxt_addr[2] .shared_arith = "off";

dffeas \int_nxt_addr_reg[2] (
	.clk(clk_clk),
	.d(\nxt_addr[2]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[2]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~1 (
	.dataa(!h2f_ARADDR_2),
	.datab(!sink0_data[69]),
	.datac(!\new_burst_reg~q ),
	.datad(!\int_nxt_addr_reg[2]~q ),
	.datae(!\in_burstwrap_reg[2]~q ),
	.dataf(!\Add0~5_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~1 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~1 .lut_mask = 64'h01F101F101F1F1F1;
defparam \d0_int_nxt_addr[2]~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_address_alignment_4 (
	new_burst_reg,
	src_payload,
	in_size_reg_0,
	src_payload1,
	in_size_reg_2,
	src_payload2,
	in_size_reg_1,
	LessThan0,
	LessThan01)/* synthesis synthesis_greybox=0 */;
input 	new_burst_reg;
input 	src_payload;
input 	in_size_reg_0;
input 	src_payload1;
input 	in_size_reg_2;
input 	src_payload2;
input 	in_size_reg_1;
output 	LessThan0;
output 	LessThan01;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!new_burst_reg),
	.datab(!src_payload1),
	.datac(!in_size_reg_2),
	.datad(!src_payload2),
	.datae(!in_size_reg_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan0),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'hE4A04400E4A04400;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~1 (
	.dataa(!new_burst_reg),
	.datab(!src_payload),
	.datac(!in_size_reg_0),
	.datad(!LessThan0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan01),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~1 .extended_lut = "off";
defparam \LessThan0~1 .lut_mask = 64'h00E400E400E400E4;
defparam \LessThan0~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_burst_adapter_4 (
	h2f_ARADDR_0,
	h2f_ARADDR_1,
	h2f_ARADDR_2,
	h2f_ARADDR_3,
	h2f_ARBURST_0,
	h2f_ARBURST_1,
	h2f_ARID_0,
	h2f_ARID_1,
	h2f_ARID_2,
	h2f_ARID_3,
	h2f_ARID_4,
	h2f_ARID_5,
	h2f_ARID_6,
	h2f_ARID_7,
	h2f_ARID_8,
	h2f_ARID_9,
	h2f_ARID_10,
	h2f_ARID_11,
	h2f_ARLEN_0,
	Add5,
	Add51,
	in_ready_hold,
	in_data_reg_69,
	stateST_COMP_TRANS,
	mem_used_1,
	in_narrow_reg,
	cp_ready,
	nxt_in_ready,
	out_valid_reg,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready1,
	saved_grant_1,
	altera_reset_synchronizer_int_chain_out,
	Decoder1,
	Add2,
	Add21,
	Add22,
	Add23,
	nxt_in_ready2,
	src_valid,
	nxt_out_eop,
	out_byte_cnt_reg_2,
	cp_ready1,
	out_uncomp_byte_cnt_reg_6,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	Selector10,
	Selector101,
	Selector11,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	Selector12,
	src_payload,
	src_payload1,
	src_payload2,
	Selector13,
	nxt_out_burstwrap_1,
	nxt_addr_2,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARADDR_0;
input 	h2f_ARADDR_1;
input 	h2f_ARADDR_2;
input 	h2f_ARADDR_3;
input 	h2f_ARBURST_0;
input 	h2f_ARBURST_1;
input 	h2f_ARID_0;
input 	h2f_ARID_1;
input 	h2f_ARID_2;
input 	h2f_ARID_3;
input 	h2f_ARID_4;
input 	h2f_ARID_5;
input 	h2f_ARID_6;
input 	h2f_ARID_7;
input 	h2f_ARID_8;
input 	h2f_ARID_9;
input 	h2f_ARID_10;
input 	h2f_ARID_11;
input 	h2f_ARLEN_0;
input 	Add5;
input 	Add51;
input 	in_ready_hold;
output 	in_data_reg_69;
output 	stateST_COMP_TRANS;
input 	mem_used_1;
output 	in_narrow_reg;
input 	cp_ready;
output 	nxt_in_ready;
output 	out_valid_reg;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready1;
input 	saved_grant_1;
input 	altera_reset_synchronizer_int_chain_out;
input 	Decoder1;
input 	Add2;
input 	Add21;
input 	Add22;
input 	Add23;
output 	nxt_in_ready2;
input 	src_valid;
output 	nxt_out_eop;
output 	out_byte_cnt_reg_2;
input 	cp_ready1;
output 	out_uncomp_byte_cnt_reg_6;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	in_data_reg_105;
output 	in_data_reg_106;
output 	in_data_reg_107;
output 	in_data_reg_108;
output 	in_data_reg_109;
output 	in_data_reg_110;
output 	in_data_reg_111;
output 	in_data_reg_112;
output 	in_data_reg_113;
output 	in_data_reg_114;
output 	in_data_reg_115;
output 	in_data_reg_116;
input 	Selector10;
input 	Selector101;
input 	Selector11;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
input 	Selector12;
input 	src_payload;
input 	src_payload1;
input 	src_payload2;
input 	Selector13;
input 	nxt_out_burstwrap_1;
input 	nxt_addr_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



spw_babasu_altera_merlin_burst_adapter_13_1_4 \altera_merlin_burst_adapter_13_1.burst_adapter (
	.h2f_ARADDR_0(h2f_ARADDR_0),
	.h2f_ARADDR_1(h2f_ARADDR_1),
	.h2f_ARADDR_2(h2f_ARADDR_2),
	.h2f_ARADDR_3(h2f_ARADDR_3),
	.h2f_ARBURST_0(h2f_ARBURST_0),
	.h2f_ARBURST_1(h2f_ARBURST_1),
	.sink0_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,h2f_ARID_11,h2f_ARID_10,h2f_ARID_9,h2f_ARID_8,h2f_ARID_7,h2f_ARID_6,h2f_ARID_5,h2f_ARID_4,h2f_ARID_3,h2f_ARID_2,h2f_ARID_1,h2f_ARID_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_payload1,src_payload2,src_payload,gnd,gnd,gnd,
Selector101,Selector11,Selector12,Selector13,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,saved_grant_1,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.h2f_ARLEN_0(h2f_ARLEN_0),
	.Add5(Add5),
	.Add51(Add51),
	.in_ready_hold(in_ready_hold),
	.in_data_reg_69(in_data_reg_69),
	.stateST_COMP_TRANS(stateST_COMP_TRANS),
	.mem_used_1(mem_used_1),
	.in_narrow_reg1(in_narrow_reg),
	.cp_ready(cp_ready),
	.nxt_in_ready(nxt_in_ready),
	.out_valid_reg1(out_valid_reg),
	.stateST_UNCOMP_WR_SUBBURST(stateST_UNCOMP_WR_SUBBURST),
	.nxt_in_ready1(nxt_in_ready1),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.Decoder1(Decoder1),
	.Add2(Add2),
	.Add21(Add21),
	.Add22(Add22),
	.Add23(Add23),
	.nxt_in_ready2(nxt_in_ready2),
	.src_valid(src_valid),
	.nxt_out_eop(nxt_out_eop),
	.out_byte_cnt_reg_2(out_byte_cnt_reg_2),
	.cp_ready1(cp_ready1),
	.out_uncomp_byte_cnt_reg_6(out_uncomp_byte_cnt_reg_6),
	.out_uncomp_byte_cnt_reg_5(out_uncomp_byte_cnt_reg_5),
	.out_uncomp_byte_cnt_reg_4(out_uncomp_byte_cnt_reg_4),
	.out_uncomp_byte_cnt_reg_3(out_uncomp_byte_cnt_reg_3),
	.out_uncomp_byte_cnt_reg_2(out_uncomp_byte_cnt_reg_2),
	.in_data_reg_105(in_data_reg_105),
	.in_data_reg_106(in_data_reg_106),
	.in_data_reg_107(in_data_reg_107),
	.in_data_reg_108(in_data_reg_108),
	.in_data_reg_109(in_data_reg_109),
	.in_data_reg_110(in_data_reg_110),
	.in_data_reg_111(in_data_reg_111),
	.in_data_reg_112(in_data_reg_112),
	.in_data_reg_113(in_data_reg_113),
	.in_data_reg_114(in_data_reg_114),
	.in_data_reg_115(in_data_reg_115),
	.in_data_reg_116(in_data_reg_116),
	.Selector10(Selector10),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_3),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_2),
	.nxt_out_burstwrap_1(nxt_out_burstwrap_1),
	.nxt_addr_2(nxt_addr_2),
	.clk_clk(clk_clk));

endmodule

module spw_babasu_altera_merlin_burst_adapter_13_1_4 (
	h2f_ARADDR_0,
	h2f_ARADDR_1,
	h2f_ARADDR_2,
	h2f_ARADDR_3,
	h2f_ARBURST_0,
	h2f_ARBURST_1,
	sink0_data,
	h2f_ARLEN_0,
	Add5,
	Add51,
	in_ready_hold,
	in_data_reg_69,
	stateST_COMP_TRANS,
	mem_used_1,
	in_narrow_reg1,
	cp_ready,
	nxt_in_ready,
	out_valid_reg1,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready1,
	altera_reset_synchronizer_int_chain_out,
	Decoder1,
	Add2,
	Add21,
	Add22,
	Add23,
	nxt_in_ready2,
	src_valid,
	nxt_out_eop,
	out_byte_cnt_reg_2,
	cp_ready1,
	out_uncomp_byte_cnt_reg_6,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	Selector10,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	nxt_out_burstwrap_1,
	nxt_addr_2,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARADDR_0;
input 	h2f_ARADDR_1;
input 	h2f_ARADDR_2;
input 	h2f_ARADDR_3;
input 	h2f_ARBURST_0;
input 	h2f_ARBURST_1;
input 	[128:0] sink0_data;
input 	h2f_ARLEN_0;
input 	Add5;
input 	Add51;
input 	in_ready_hold;
output 	in_data_reg_69;
output 	stateST_COMP_TRANS;
input 	mem_used_1;
output 	in_narrow_reg1;
input 	cp_ready;
output 	nxt_in_ready;
output 	out_valid_reg1;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready1;
input 	altera_reset_synchronizer_int_chain_out;
input 	Decoder1;
input 	Add2;
input 	Add21;
input 	Add22;
input 	Add23;
output 	nxt_in_ready2;
input 	src_valid;
output 	nxt_out_eop;
output 	out_byte_cnt_reg_2;
input 	cp_ready1;
output 	out_uncomp_byte_cnt_reg_6;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	in_data_reg_105;
output 	in_data_reg_106;
output 	in_data_reg_107;
output 	in_data_reg_108;
output 	in_data_reg_109;
output 	in_data_reg_110;
output 	in_data_reg_111;
output 	in_data_reg_112;
output 	in_data_reg_113;
output 	in_data_reg_114;
output 	in_data_reg_115;
output 	in_data_reg_116;
input 	Selector10;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
input 	nxt_out_burstwrap_1;
input 	nxt_addr_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \align_address_to_size|LessThan0~0_combout ;
wire \align_address_to_size|LessThan0~1_combout ;
wire \NON_PIPELINED_INPUTS.load_next_cmd~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt~0_combout ;
wire \Add4~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt[6]~1_combout ;
wire \nxt_uncomp_subburst_byte_cnt[5]~2_combout ;
wire \nxt_uncomp_subburst_byte_cnt[4]~3_combout ;
wire \nxt_uncomp_subburst_byte_cnt[3]~4_combout ;
wire \nxt_uncomp_subburst_byte_cnt[2]~5_combout ;
wire \WideNor1~combout ;
wire \Selector2~1_combout ;
wire \load_next_out_cmd~combout ;
wire \state.ST_UNCOMP_TRANS~q ;
wire \Selector2~0_combout ;
wire \Selector0~0_combout ;
wire \state.ST_IDLE~q ;
wire \Selector1~0_combout ;
wire \Selector1~1_combout ;
wire \int_bytes_remaining_reg[5]~q ;
wire \d0_int_bytes_remaining[2]~4_combout ;
wire \int_bytes_remaining_reg[2]~q ;
wire \d0_int_bytes_remaining[3]~3_combout ;
wire \int_bytes_remaining_reg[3]~q ;
wire \Add1~1_combout ;
wire \d0_int_bytes_remaining[4]~2_combout ;
wire \int_bytes_remaining_reg[4]~q ;
wire \Add1~0_combout ;
wire \d0_int_bytes_remaining[5]~0_combout ;
wire \int_bytes_remaining_reg[6]~q ;
wire \d0_int_bytes_remaining[6]~1_combout ;
wire \new_burst_reg~0_combout ;
wire \new_burst_reg~q ;
wire \in_bytecount_reg_zero~0_combout ;
wire \in_bytecount_reg_zero~q ;
wire \nxt_out_valid~0_combout ;
wire \nxt_out_valid~1_combout ;
wire \Selector3~0_combout ;
wire \in_burstwrap_reg[3]~q ;
wire \nxt_addr[3]~0_combout ;
wire \nxt_addr[3]~combout ;
wire \int_nxt_addr_reg[3]~q ;
wire \in_size_reg[0]~q ;
wire \in_size_reg[2]~q ;
wire \in_size_reg[1]~q ;
wire \ShiftLeft0~0_combout ;
wire \ShiftLeft0~1_combout ;
wire \int_byte_cnt_narrow_reg[3]~q ;
wire \ShiftLeft0~2_combout ;
wire \int_byte_cnt_narrow_reg[2]~q ;
wire \in_burstwrap_reg[1]~q ;
wire \nxt_addr[1]~combout ;
wire \int_nxt_addr_reg[1]~q ;
wire \ShiftLeft0~3_combout ;
wire \int_byte_cnt_narrow_reg[1]~q ;
wire \int_byte_cnt_narrow_reg[0]~q ;
wire \Add0~13_sumout ;
wire \in_burstwrap_reg[0]~q ;
wire \nxt_addr[0]~combout ;
wire \int_nxt_addr_reg[0]~q ;
wire \d0_int_nxt_addr[0]~2_combout ;
wire \d0_int_nxt_addr[0]~3_combout ;
wire \int_nxt_addr_reg_dly[0]~q ;
wire \Add0~14 ;
wire \Add0~9_sumout ;
wire \d0_int_nxt_addr[1]~4_combout ;
wire \int_nxt_addr_reg_dly[1]~q ;
wire \Add0~10 ;
wire \Add0~6 ;
wire \Add0~1_sumout ;
wire \d0_int_nxt_addr[3]~0_combout ;
wire \in_burstwrap_reg[2]~q ;
wire \nxt_addr[2]~1_combout ;
wire \nxt_addr[2]~combout ;
wire \int_nxt_addr_reg[2]~q ;
wire \Add0~5_sumout ;
wire \d0_int_nxt_addr[2]~1_combout ;


spw_babasu_altera_merlin_address_alignment_5 align_address_to_size(
	.new_burst_reg(\new_burst_reg~q ),
	.src_payload(sink0_data[86]),
	.in_size_reg_0(\in_size_reg[0]~q ),
	.src_payload1(sink0_data[88]),
	.in_size_reg_2(\in_size_reg[2]~q ),
	.src_payload2(sink0_data[87]),
	.in_size_reg_1(\in_size_reg[1]~q ),
	.LessThan0(\align_address_to_size|LessThan0~0_combout ),
	.LessThan01(\align_address_to_size|LessThan0~1_combout ));

dffeas \in_data_reg[69] (
	.clk(clk_clk),
	.d(sink0_data[69]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_69),
	.prn(vcc));
defparam \in_data_reg[69] .is_wysiwyg = "true";
defparam \in_data_reg[69] .power_up = "low";

dffeas \state.ST_COMP_TRANS (
	.clk(clk_clk),
	.d(\Selector1~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_COMP_TRANS),
	.prn(vcc));
defparam \state.ST_COMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_COMP_TRANS .power_up = "low";

dffeas in_narrow_reg(
	.clk(clk_clk),
	.d(Decoder1),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_narrow_reg1),
	.prn(vcc));
defparam in_narrow_reg.is_wysiwyg = "true";
defparam in_narrow_reg.power_up = "low";

cyclonev_lcell_comb \nxt_in_ready~0 (
	.dataa(gnd),
	.datab(!stateST_COMP_TRANS),
	.datac(!\new_burst_reg~q ),
	.datad(!mem_used_1),
	.datae(!cp_ready),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~0 .extended_lut = "off";
defparam \nxt_in_ready~0 .lut_mask = 64'h0000030000000300;
defparam \nxt_in_ready~0 .shared_arith = "off";

dffeas out_valid_reg(
	.clk(clk_clk),
	.d(\nxt_out_valid~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_valid_reg1),
	.prn(vcc));
defparam out_valid_reg.is_wysiwyg = "true";
defparam out_valid_reg.power_up = "low";

dffeas \state.ST_UNCOMP_WR_SUBBURST (
	.clk(clk_clk),
	.d(\Selector3~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_UNCOMP_WR_SUBBURST),
	.prn(vcc));
defparam \state.ST_UNCOMP_WR_SUBBURST .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_WR_SUBBURST .power_up = "low";

cyclonev_lcell_comb \nxt_in_ready~1 (
	.dataa(!in_ready_hold),
	.datab(!stateST_COMP_TRANS),
	.datac(!mem_used_1),
	.datad(!cp_ready),
	.datae(!out_valid_reg1),
	.dataf(!\Selector2~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~1 .extended_lut = "off";
defparam \nxt_in_ready~1 .lut_mask = 64'h0000FF3F8888BBBB;
defparam \nxt_in_ready~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_in_ready~2 (
	.dataa(!nxt_in_ready),
	.datab(!nxt_in_ready1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready2),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~2 .extended_lut = "off";
defparam \nxt_in_ready~2 .lut_mask = 64'h2222222222222222;
defparam \nxt_in_ready~2 .shared_arith = "off";

cyclonev_lcell_comb \nxt_out_eop~0 (
	.dataa(!in_data_reg_69),
	.datab(!stateST_COMP_TRANS),
	.datac(!\new_burst_reg~q ),
	.datad(!mem_used_1),
	.datae(!cp_ready),
	.dataf(!\in_bytecount_reg_zero~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_out_eop),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_eop~0 .extended_lut = "off";
defparam \nxt_out_eop~0 .lut_mask = 64'h4444474477774777;
defparam \nxt_out_eop~0 .shared_arith = "off";

dffeas \out_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[6] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[6]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_6),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[6] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[6] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[5] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[5]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_5),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[5] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[5] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[4] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[4]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_4),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[4] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[4] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[3] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[3]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_3),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[3] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[3] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[2]~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[2] .power_up = "low";

dffeas \in_data_reg[105] (
	.clk(clk_clk),
	.d(sink0_data[105]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_105),
	.prn(vcc));
defparam \in_data_reg[105] .is_wysiwyg = "true";
defparam \in_data_reg[105] .power_up = "low";

dffeas \in_data_reg[106] (
	.clk(clk_clk),
	.d(sink0_data[106]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_106),
	.prn(vcc));
defparam \in_data_reg[106] .is_wysiwyg = "true";
defparam \in_data_reg[106] .power_up = "low";

dffeas \in_data_reg[107] (
	.clk(clk_clk),
	.d(sink0_data[107]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_107),
	.prn(vcc));
defparam \in_data_reg[107] .is_wysiwyg = "true";
defparam \in_data_reg[107] .power_up = "low";

dffeas \in_data_reg[108] (
	.clk(clk_clk),
	.d(sink0_data[108]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_108),
	.prn(vcc));
defparam \in_data_reg[108] .is_wysiwyg = "true";
defparam \in_data_reg[108] .power_up = "low";

dffeas \in_data_reg[109] (
	.clk(clk_clk),
	.d(sink0_data[109]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_109),
	.prn(vcc));
defparam \in_data_reg[109] .is_wysiwyg = "true";
defparam \in_data_reg[109] .power_up = "low";

dffeas \in_data_reg[110] (
	.clk(clk_clk),
	.d(sink0_data[110]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_110),
	.prn(vcc));
defparam \in_data_reg[110] .is_wysiwyg = "true";
defparam \in_data_reg[110] .power_up = "low";

dffeas \in_data_reg[111] (
	.clk(clk_clk),
	.d(sink0_data[111]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_111),
	.prn(vcc));
defparam \in_data_reg[111] .is_wysiwyg = "true";
defparam \in_data_reg[111] .power_up = "low";

dffeas \in_data_reg[112] (
	.clk(clk_clk),
	.d(sink0_data[112]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_112),
	.prn(vcc));
defparam \in_data_reg[112] .is_wysiwyg = "true";
defparam \in_data_reg[112] .power_up = "low";

dffeas \in_data_reg[113] (
	.clk(clk_clk),
	.d(sink0_data[113]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_113),
	.prn(vcc));
defparam \in_data_reg[113] .is_wysiwyg = "true";
defparam \in_data_reg[113] .power_up = "low";

dffeas \in_data_reg[114] (
	.clk(clk_clk),
	.d(sink0_data[114]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_114),
	.prn(vcc));
defparam \in_data_reg[114] .is_wysiwyg = "true";
defparam \in_data_reg[114] .power_up = "low";

dffeas \in_data_reg[115] (
	.clk(clk_clk),
	.d(sink0_data[115]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_115),
	.prn(vcc));
defparam \in_data_reg[115] .is_wysiwyg = "true";
defparam \in_data_reg[115] .power_up = "low";

dffeas \in_data_reg[116] (
	.clk(clk_clk),
	.d(sink0_data[116]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_116),
	.prn(vcc));
defparam \in_data_reg[116] .is_wysiwyg = "true";
defparam \in_data_reg[116] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[3] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[3]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_3),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[3] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[2] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[2]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_2),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[2] .power_up = "low";

cyclonev_lcell_comb \NON_PIPELINED_INPUTS.load_next_cmd~0 (
	.dataa(!in_ready_hold),
	.datab(!nxt_in_ready2),
	.datac(!src_valid),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \NON_PIPELINED_INPUTS.load_next_cmd~0 .extended_lut = "off";
defparam \NON_PIPELINED_INPUTS.load_next_cmd~0 .lut_mask = 64'h0404040404040404;
defparam \NON_PIPELINED_INPUTS.load_next_cmd~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt~0 (
	.dataa(!mem_used_1),
	.datab(!cp_ready),
	.datac(!out_valid_reg1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt~0 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt~0 .lut_mask = 64'h0202020202020202;
defparam \nxt_uncomp_subburst_byte_cnt~0 .shared_arith = "off";

cyclonev_lcell_comb \Add4~0 (
	.dataa(!out_uncomp_byte_cnt_reg_4),
	.datab(!out_uncomp_byte_cnt_reg_3),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add4~0 .extended_lut = "off";
defparam \Add4~0 .lut_mask = 64'h0800080008000800;
defparam \Add4~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[6]~1 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_6),
	.datad(!out_uncomp_byte_cnt_reg_5),
	.datae(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.dataf(!\Add4~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[6]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[6]~1 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[6]~1 .lut_mask = 64'h0F0F4E4EA50FE44E;
defparam \nxt_uncomp_subburst_byte_cnt[6]~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[5]~2 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!\Add4~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[5]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[5]~2 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[5]~2 .lut_mask = 64'h0F4EA5E40F4EA5E4;
defparam \nxt_uncomp_subburst_byte_cnt[5]~2 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[4]~3 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!out_uncomp_byte_cnt_reg_3),
	.datae(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.dataf(!out_uncomp_byte_cnt_reg_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[4]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[4]~3 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[4]~3 .lut_mask = 64'h0F0FE44E0F0F4E4E;
defparam \nxt_uncomp_subburst_byte_cnt[4]~3 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[3]~4 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!out_uncomp_byte_cnt_reg_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[3]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[3]~4 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[3]~4 .lut_mask = 64'h0FE40F4E0FE40F4E;
defparam \nxt_uncomp_subburst_byte_cnt[3]~4 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[2]~5 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[2]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[2]~5 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[2]~5 .lut_mask = 64'h0EF40EF40EF40EF4;
defparam \nxt_uncomp_subburst_byte_cnt[2]~5 .shared_arith = "off";

cyclonev_lcell_comb WideNor1(
	.dataa(!\nxt_uncomp_subburst_byte_cnt[6]~1_combout ),
	.datab(!\nxt_uncomp_subburst_byte_cnt[5]~2_combout ),
	.datac(!\nxt_uncomp_subburst_byte_cnt[4]~3_combout ),
	.datad(!\nxt_uncomp_subburst_byte_cnt[3]~4_combout ),
	.datae(!\nxt_uncomp_subburst_byte_cnt[2]~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideNor1.extended_lut = "off";
defparam WideNor1.lut_mask = 64'h8000000080000000;
defparam WideNor1.shared_arith = "off";

cyclonev_lcell_comb \Selector2~1 (
	.dataa(!nxt_out_eop),
	.datab(!\Selector2~0_combout ),
	.datac(!\WideNor1~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~1 .extended_lut = "off";
defparam \Selector2~1 .lut_mask = 64'h0808080808080808;
defparam \Selector2~1 .shared_arith = "off";

cyclonev_lcell_comb load_next_out_cmd(
	.dataa(!mem_used_1),
	.datab(!cp_ready),
	.datac(!out_valid_reg1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\load_next_out_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam load_next_out_cmd.extended_lut = "off";
defparam load_next_out_cmd.lut_mask = 64'hF2F2F2F2F2F2F2F2;
defparam load_next_out_cmd.shared_arith = "off";

dffeas \state.ST_UNCOMP_TRANS (
	.clk(clk_clk),
	.d(\Selector2~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_UNCOMP_TRANS~q ),
	.prn(vcc));
defparam \state.ST_UNCOMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_TRANS .power_up = "low";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'h8888888888888888;
defparam \Selector2~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!in_ready_hold),
	.datab(!nxt_out_eop),
	.datac(!src_valid),
	.datad(!\state.ST_IDLE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'h05CD05CD05CD05CD;
defparam \Selector0~0 .shared_arith = "off";

dffeas \state.ST_IDLE (
	.clk(clk_clk),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_IDLE~q ),
	.prn(vcc));
defparam \state.ST_IDLE .is_wysiwyg = "true";
defparam \state.ST_IDLE .power_up = "low";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!sink0_data[69]),
	.datab(!nxt_out_eop),
	.datac(!\Selector2~0_combout ),
	.datad(!\state.ST_IDLE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'h5510551055105510;
defparam \Selector1~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~1 (
	.dataa(!in_ready_hold),
	.datab(!stateST_COMP_TRANS),
	.datac(!nxt_out_eop),
	.datad(!src_valid),
	.datae(!\Selector1~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~1 .extended_lut = "off";
defparam \Selector1~1 .lut_mask = 64'h3031307530313075;
defparam \Selector1~1 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[5] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[5]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[5]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[5] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[5] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[2]~4 (
	.dataa(!h2f_ARLEN_0),
	.datab(!sink0_data[69]),
	.datac(!\new_burst_reg~q ),
	.datad(!out_byte_cnt_reg_2),
	.datae(!\int_bytes_remaining_reg[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[2]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[2]~4 .extended_lut = "off";
defparam \d0_int_bytes_remaining[2]~4 .lut_mask = 64'h02F2F20202F2F202;
defparam \d0_int_bytes_remaining[2]~4 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[2] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[2]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[2]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[2] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[3]~3 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!Add2),
	.datad(!\int_bytes_remaining_reg[3]~q ),
	.datae(!out_byte_cnt_reg_2),
	.dataf(!\int_bytes_remaining_reg[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[3]~3 .extended_lut = "off";
defparam \d0_int_bytes_remaining[3]~3 .lut_mask = 64'h01CDCD0101CD01CD;
defparam \d0_int_bytes_remaining[3]~3 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[3] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[3]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[3]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[3] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[3] .power_up = "low";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!\int_bytes_remaining_reg[4]~q ),
	.datab(!\int_bytes_remaining_reg[3]~q ),
	.datac(!out_byte_cnt_reg_2),
	.datad(!\int_bytes_remaining_reg[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'hA6AAA6AAA6AAA6AA;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[4]~2 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!Add21),
	.datad(!\Add1~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[4]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[4]~2 .extended_lut = "off";
defparam \d0_int_bytes_remaining[4]~2 .lut_mask = 64'hCD01CD01CD01CD01;
defparam \d0_int_bytes_remaining[4]~2 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[4] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[4]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[4]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[4] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[4] .power_up = "low";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!\int_bytes_remaining_reg[4]~q ),
	.datab(!\int_bytes_remaining_reg[3]~q ),
	.datac(!out_byte_cnt_reg_2),
	.datad(!\int_bytes_remaining_reg[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h0800080008000800;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[5]~0 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!Add22),
	.datad(!\int_bytes_remaining_reg[5]~q ),
	.datae(!\Add1~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[5]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[5]~0 .extended_lut = "off";
defparam \d0_int_bytes_remaining[5]~0 .lut_mask = 64'h01CDCD0101CDCD01;
defparam \d0_int_bytes_remaining[5]~0 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[6] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[6]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[6]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[6] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[6] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[6]~1 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!Add23),
	.datad(!\int_bytes_remaining_reg[5]~q ),
	.datae(!\Add1~0_combout ),
	.dataf(!\int_bytes_remaining_reg[6]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[6]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[6]~1 .extended_lut = "off";
defparam \d0_int_bytes_remaining[6]~1 .lut_mask = 64'h0101CD01CDCD01CD;
defparam \d0_int_bytes_remaining[6]~1 .shared_arith = "off";

cyclonev_lcell_comb \new_burst_reg~0 (
	.dataa(!\Selector1~1_combout ),
	.datab(!\d0_int_bytes_remaining[5]~0_combout ),
	.datac(!\d0_int_bytes_remaining[6]~1_combout ),
	.datad(!\d0_int_bytes_remaining[4]~2_combout ),
	.datae(!\d0_int_bytes_remaining[3]~3_combout ),
	.dataf(!\d0_int_bytes_remaining[2]~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\new_burst_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \new_burst_reg~0 .extended_lut = "off";
defparam \new_burst_reg~0 .lut_mask = 64'hAAAAAAAAEAAAAAAA;
defparam \new_burst_reg~0 .shared_arith = "off";

dffeas new_burst_reg(
	.clk(clk_clk),
	.d(\new_burst_reg~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\new_burst_reg~q ),
	.prn(vcc));
defparam new_burst_reg.is_wysiwyg = "true";
defparam new_burst_reg.power_up = "low";

cyclonev_lcell_comb \in_bytecount_reg_zero~0 (
	.dataa(!sink0_data[69]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\in_bytecount_reg_zero~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \in_bytecount_reg_zero~0 .extended_lut = "off";
defparam \in_bytecount_reg_zero~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \in_bytecount_reg_zero~0 .shared_arith = "off";

dffeas in_bytecount_reg_zero(
	.clk(clk_clk),
	.d(\in_bytecount_reg_zero~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_bytecount_reg_zero~q ),
	.prn(vcc));
defparam in_bytecount_reg_zero.is_wysiwyg = "true";
defparam in_bytecount_reg_zero.power_up = "low";

cyclonev_lcell_comb \nxt_out_valid~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!mem_used_1),
	.datac(!\in_bytecount_reg_zero~q ),
	.datad(!cp_ready1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_valid~0 .extended_lut = "off";
defparam \nxt_out_valid~0 .lut_mask = 64'hF0B8F0B8F0B8F0B8;
defparam \nxt_out_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_out_valid~1 (
	.dataa(!in_ready_hold),
	.datab(!stateST_COMP_TRANS),
	.datac(!src_valid),
	.datad(!\nxt_out_valid~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_valid~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_valid~1 .extended_lut = "off";
defparam \nxt_out_valid~1 .lut_mask = 64'h0537053705370537;
defparam \nxt_out_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~0 (
	.dataa(!nxt_out_eop),
	.datab(!\Selector2~0_combout ),
	.datac(!\WideNor1~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'h8080808080808080;
defparam \Selector3~0 .shared_arith = "off";

dffeas \in_burstwrap_reg[3] (
	.clk(clk_clk),
	.d(sink0_data[82]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_burstwrap_reg[3]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[3] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[3] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[3]~0 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!\in_burstwrap_reg[3]~q ),
	.datad(!\d0_int_nxt_addr[3]~0_combout ),
	.datae(!h2f_ARBURST_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[3]~0 .extended_lut = "off";
defparam \nxt_addr[3]~0 .lut_mask = 64'h00F300E200F300E2;
defparam \nxt_addr[3]~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_addr[3] (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!h2f_ARBURST_1),
	.datad(!Add5),
	.datae(!Selector10),
	.dataf(!\nxt_addr[3]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[3] .extended_lut = "off";
defparam \nxt_addr[3] .lut_mask = 64'h00000000FEEEFFEF;
defparam \nxt_addr[3] .shared_arith = "off";

dffeas \int_nxt_addr_reg[3] (
	.clk(clk_clk),
	.d(\nxt_addr[3]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[3]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[3] .power_up = "low";

dffeas \in_size_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[86]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_size_reg[0]~q ),
	.prn(vcc));
defparam \in_size_reg[0] .is_wysiwyg = "true";
defparam \in_size_reg[0] .power_up = "low";

dffeas \in_size_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[88]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_size_reg[2]~q ),
	.prn(vcc));
defparam \in_size_reg[2] .is_wysiwyg = "true";
defparam \in_size_reg[2] .power_up = "low";

dffeas \in_size_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[87]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_size_reg[1]~q ),
	.prn(vcc));
defparam \in_size_reg[1] .is_wysiwyg = "true";
defparam \in_size_reg[1] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[88]),
	.datac(!\in_size_reg[2]~q ),
	.datad(!sink0_data[87]),
	.datae(!\in_size_reg[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~0 .extended_lut = "off";
defparam \ShiftLeft0~0 .lut_mask = 64'h0044A0E40044A0E4;
defparam \ShiftLeft0~0 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~1 .extended_lut = "off";
defparam \ShiftLeft0~1 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~1 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[3] (
	.clk(clk_clk),
	.d(\ShiftLeft0~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[3]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[3] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[3] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~2 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~2 .extended_lut = "off";
defparam \ShiftLeft0~2 .lut_mask = 64'h00E400E400E400E4;
defparam \ShiftLeft0~2 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[2] (
	.clk(clk_clk),
	.d(\ShiftLeft0~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[2]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[2] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[2] .power_up = "low";

dffeas \in_burstwrap_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[80]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_burstwrap_reg[1]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[1] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[1] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[1] (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!\in_burstwrap_reg[1]~q ),
	.datad(!\d0_int_nxt_addr[1]~4_combout ),
	.datae(!nxt_out_burstwrap_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[1] .extended_lut = "off";
defparam \nxt_addr[1] .lut_mask = 64'h00E200F300E200F3;
defparam \nxt_addr[1] .shared_arith = "off";

dffeas \int_nxt_addr_reg[1] (
	.clk(clk_clk),
	.d(\nxt_addr[1]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[1] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\align_address_to_size|LessThan0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~3 .extended_lut = "off";
defparam \ShiftLeft0~3 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~3 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[1] (
	.clk(clk_clk),
	.d(\ShiftLeft0~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[1]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[1] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[1] .power_up = "low";

dffeas \int_byte_cnt_narrow_reg[0] (
	.clk(clk_clk),
	.d(\align_address_to_size|LessThan0~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[0]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[0] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[0] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[0]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \in_burstwrap_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[79]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_burstwrap_reg[0]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[0] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[0] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[0] (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!sink0_data[79]),
	.datad(!\in_burstwrap_reg[0]~q ),
	.datae(!\d0_int_nxt_addr[0]~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[0] .extended_lut = "off";
defparam \nxt_addr[0] .lut_mask = 64'h0000FE320000FE32;
defparam \nxt_addr[0] .shared_arith = "off";

dffeas \int_nxt_addr_reg[0] (
	.clk(clk_clk),
	.d(\nxt_addr[0]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[0] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~2 (
	.dataa(!\Add0~13_sumout ),
	.datab(!\int_nxt_addr_reg[0]~q ),
	.datac(!\in_burstwrap_reg[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~2 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~2 .lut_mask = 64'hC8C8C8C8C8C8C8C8;
defparam \d0_int_nxt_addr[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~3 (
	.dataa(!h2f_ARADDR_0),
	.datab(!sink0_data[69]),
	.datac(!\new_burst_reg~q ),
	.datad(!\align_address_to_size|LessThan0~1_combout ),
	.datae(!\d0_int_nxt_addr[0]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~3 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~3 .lut_mask = 64'hF0F10001F0F10001;
defparam \d0_int_nxt_addr[0]~3 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[0] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[0]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[0] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[1]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[1]~q ),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~4 (
	.dataa(!\int_nxt_addr_reg[1]~q ),
	.datab(!\Add0~9_sumout ),
	.datac(!sink0_data[69]),
	.datad(!Decoder1),
	.datae(!\new_burst_reg~q ),
	.dataf(!h2f_ARADDR_1),
	.datag(!\in_burstwrap_reg[1]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~4 .extended_lut = "on";
defparam \d0_int_nxt_addr[1]~4 .lut_mask = 64'h575700005757000F;
defparam \d0_int_nxt_addr[1]~4 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[1] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[1]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[1] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_2),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[2]~q ),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[3]~q ),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~0 (
	.dataa(!h2f_ARADDR_3),
	.datab(!sink0_data[69]),
	.datac(!\new_burst_reg~q ),
	.datad(!\int_nxt_addr_reg[3]~q ),
	.datae(!\in_burstwrap_reg[3]~q ),
	.dataf(!\Add0~1_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~0 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~0 .lut_mask = 64'h01F101F101F1F1F1;
defparam \d0_int_nxt_addr[3]~0 .shared_arith = "off";

dffeas \in_burstwrap_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[81]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_burstwrap_reg[2]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[2] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[2] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[2]~1 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!\in_burstwrap_reg[2]~q ),
	.datad(!\d0_int_nxt_addr[2]~1_combout ),
	.datae(!h2f_ARBURST_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[2]~1 .extended_lut = "off";
defparam \nxt_addr[2]~1 .lut_mask = 64'h00F300E200F300E2;
defparam \nxt_addr[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_addr[2] (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!h2f_ARBURST_1),
	.datad(!Add51),
	.datae(!\nxt_addr[2]~1_combout ),
	.dataf(!nxt_addr_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[2] .extended_lut = "off";
defparam \nxt_addr[2] .lut_mask = 64'h0000FEEE0000FFEF;
defparam \nxt_addr[2] .shared_arith = "off";

dffeas \int_nxt_addr_reg[2] (
	.clk(clk_clk),
	.d(\nxt_addr[2]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[2]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~1 (
	.dataa(!h2f_ARADDR_2),
	.datab(!sink0_data[69]),
	.datac(!\new_burst_reg~q ),
	.datad(!\int_nxt_addr_reg[2]~q ),
	.datae(!\in_burstwrap_reg[2]~q ),
	.dataf(!\Add0~5_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~1 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~1 .lut_mask = 64'h01F101F101F1F1F1;
defparam \d0_int_nxt_addr[2]~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_address_alignment_5 (
	new_burst_reg,
	src_payload,
	in_size_reg_0,
	src_payload1,
	in_size_reg_2,
	src_payload2,
	in_size_reg_1,
	LessThan0,
	LessThan01)/* synthesis synthesis_greybox=0 */;
input 	new_burst_reg;
input 	src_payload;
input 	in_size_reg_0;
input 	src_payload1;
input 	in_size_reg_2;
input 	src_payload2;
input 	in_size_reg_1;
output 	LessThan0;
output 	LessThan01;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!new_burst_reg),
	.datab(!src_payload1),
	.datac(!in_size_reg_2),
	.datad(!src_payload2),
	.datae(!in_size_reg_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan0),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'hE4A04400E4A04400;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~1 (
	.dataa(!new_burst_reg),
	.datab(!src_payload),
	.datac(!in_size_reg_0),
	.datad(!LessThan0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan01),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~1 .extended_lut = "off";
defparam \LessThan0~1 .lut_mask = 64'h00E400E400E400E4;
defparam \LessThan0~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_burst_adapter_5 (
	h2f_ARADDR_0,
	h2f_ARADDR_1,
	h2f_ARADDR_2,
	h2f_ARADDR_3,
	h2f_ARLEN_0,
	nxt_in_ready,
	in_ready_hold,
	stateST_COMP_TRANS,
	out_valid_reg,
	in_narrow_reg,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	in_data_reg_68,
	cp_ready,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready1,
	saved_grant_1,
	Equal16,
	saved_grant_0,
	altera_reset_synchronizer_int_chain_out,
	in_data_reg_0,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	Add2,
	Add21,
	Add22,
	Add23,
	nxt_out_eop,
	Equal5,
	src1_valid,
	src_valid,
	cp_ready1,
	in_data_reg_69,
	src_data_87,
	src_data_88,
	src_valid1,
	src_data_35,
	src_data_34,
	src_data_33,
	src_data_32,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_6,
	src_payload_0,
	write_cp_data_77,
	write_cp_data_78,
	write_cp_data_75,
	write_cp_data_74,
	write_cp_data_76,
	WideNor0,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	Selector3,
	Selector10,
	base_address_3,
	Selector4,
	Selector11,
	base_address_2,
	src_payload,
	src_data_82,
	src_data_81,
	src_data_105,
	src_data_106,
	src_data_107,
	src_data_108,
	src_data_109,
	src_data_110,
	src_data_111,
	src_data_112,
	src_data_113,
	src_data_114,
	src_data_115,
	src_data_116,
	src_data_86,
	Selector5,
	Selector12,
	out_data_1,
	src_data_80,
	out_data_0,
	Selector6,
	Selector13,
	src_data_79,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARADDR_0;
input 	h2f_ARADDR_1;
input 	h2f_ARADDR_2;
input 	h2f_ARADDR_3;
input 	h2f_ARLEN_0;
output 	nxt_in_ready;
input 	in_ready_hold;
output 	stateST_COMP_TRANS;
output 	out_valid_reg;
output 	in_narrow_reg;
output 	in_byteen_reg_3;
output 	in_byteen_reg_2;
output 	in_byteen_reg_1;
output 	in_byteen_reg_0;
output 	in_data_reg_68;
input 	cp_ready;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready1;
input 	saved_grant_1;
input 	Equal16;
input 	saved_grant_0;
input 	altera_reset_synchronizer_int_chain_out;
output 	in_data_reg_0;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
input 	Add2;
input 	Add21;
input 	Add22;
input 	Add23;
output 	nxt_out_eop;
input 	Equal5;
input 	src1_valid;
input 	src_valid;
input 	cp_ready1;
output 	in_data_reg_69;
input 	src_data_87;
input 	src_data_88;
input 	src_valid1;
input 	src_data_35;
input 	src_data_34;
input 	src_data_33;
input 	src_data_32;
output 	out_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_6;
input 	src_payload_0;
input 	write_cp_data_77;
input 	write_cp_data_78;
input 	write_cp_data_75;
input 	write_cp_data_74;
input 	write_cp_data_76;
input 	WideNor0;
output 	in_data_reg_105;
output 	in_data_reg_106;
output 	in_data_reg_107;
output 	in_data_reg_108;
output 	in_data_reg_109;
output 	in_data_reg_110;
output 	in_data_reg_111;
output 	in_data_reg_112;
output 	in_data_reg_113;
output 	in_data_reg_114;
output 	in_data_reg_115;
output 	in_data_reg_116;
input 	Selector3;
input 	Selector10;
input 	base_address_3;
input 	Selector4;
input 	Selector11;
input 	base_address_2;
input 	src_payload;
input 	src_data_82;
input 	src_data_81;
input 	src_data_105;
input 	src_data_106;
input 	src_data_107;
input 	src_data_108;
input 	src_data_109;
input 	src_data_110;
input 	src_data_111;
input 	src_data_112;
input 	src_data_113;
input 	src_data_114;
input 	src_data_115;
input 	src_data_116;
input 	src_data_86;
input 	Selector5;
input 	Selector12;
input 	out_data_1;
input 	src_data_80;
input 	out_data_0;
input 	Selector6;
input 	Selector13;
input 	src_data_79;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



spw_babasu_altera_merlin_burst_adapter_13_1_5 \altera_merlin_burst_adapter_13_1.burst_adapter (
	.h2f_ARADDR_0(h2f_ARADDR_0),
	.h2f_ARADDR_1(h2f_ARADDR_1),
	.h2f_ARADDR_2(h2f_ARADDR_2),
	.h2f_ARADDR_3(h2f_ARADDR_3),
	.h2f_ARLEN_0(h2f_ARLEN_0),
	.nxt_in_ready(nxt_in_ready),
	.in_ready_hold(in_ready_hold),
	.stateST_COMP_TRANS(stateST_COMP_TRANS),
	.out_valid_reg1(out_valid_reg),
	.in_narrow_reg1(in_narrow_reg),
	.in_byteen_reg_3(in_byteen_reg_3),
	.in_byteen_reg_2(in_byteen_reg_2),
	.in_byteen_reg_1(in_byteen_reg_1),
	.in_byteen_reg_0(in_byteen_reg_0),
	.in_data_reg_68(in_data_reg_68),
	.cp_ready(cp_ready),
	.stateST_UNCOMP_WR_SUBBURST(stateST_UNCOMP_WR_SUBBURST),
	.nxt_in_ready1(nxt_in_ready1),
	.sink0_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_116,src_data_115,src_data_114,src_data_113,src_data_112,src_data_111,src_data_110,src_data_109,src_data_108,src_data_107,src_data_106,src_data_105,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_88,src_data_87,
src_data_86,gnd,gnd,gnd,src_data_82,src_data_81,src_data_80,src_data_79,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,saved_grant_1,saved_grant_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_35,src_data_34,src_data_33,
src_data_32,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_payload}),
	.Equal16(Equal16),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.in_data_reg_0(in_data_reg_0),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_3),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_2),
	.Add2(Add2),
	.Add21(Add21),
	.Add22(Add22),
	.Add23(Add23),
	.nxt_out_eop(nxt_out_eop),
	.Equal5(Equal5),
	.src1_valid(src1_valid),
	.src_valid(src_valid),
	.cp_ready1(cp_ready1),
	.in_data_reg_69(in_data_reg_69),
	.src_valid1(src_valid1),
	.out_byte_cnt_reg_2(out_byte_cnt_reg_2),
	.out_uncomp_byte_cnt_reg_3(out_uncomp_byte_cnt_reg_3),
	.out_uncomp_byte_cnt_reg_2(out_uncomp_byte_cnt_reg_2),
	.out_uncomp_byte_cnt_reg_4(out_uncomp_byte_cnt_reg_4),
	.out_uncomp_byte_cnt_reg_5(out_uncomp_byte_cnt_reg_5),
	.out_uncomp_byte_cnt_reg_6(out_uncomp_byte_cnt_reg_6),
	.sink0_endofpacket(src_payload_0),
	.write_cp_data_77(write_cp_data_77),
	.write_cp_data_78(write_cp_data_78),
	.write_cp_data_75(write_cp_data_75),
	.write_cp_data_74(write_cp_data_74),
	.write_cp_data_76(write_cp_data_76),
	.WideNor0(WideNor0),
	.in_data_reg_105(in_data_reg_105),
	.in_data_reg_106(in_data_reg_106),
	.in_data_reg_107(in_data_reg_107),
	.in_data_reg_108(in_data_reg_108),
	.in_data_reg_109(in_data_reg_109),
	.in_data_reg_110(in_data_reg_110),
	.in_data_reg_111(in_data_reg_111),
	.in_data_reg_112(in_data_reg_112),
	.in_data_reg_113(in_data_reg_113),
	.in_data_reg_114(in_data_reg_114),
	.in_data_reg_115(in_data_reg_115),
	.in_data_reg_116(in_data_reg_116),
	.Selector3(Selector3),
	.Selector10(Selector10),
	.base_address_3(base_address_3),
	.Selector4(Selector4),
	.Selector11(Selector11),
	.base_address_2(base_address_2),
	.Selector5(Selector5),
	.Selector12(Selector12),
	.out_data_1(out_data_1),
	.out_data_0(out_data_0),
	.Selector6(Selector6),
	.Selector13(Selector13),
	.clk_clk(clk_clk));

endmodule

module spw_babasu_altera_merlin_burst_adapter_13_1_5 (
	h2f_ARADDR_0,
	h2f_ARADDR_1,
	h2f_ARADDR_2,
	h2f_ARADDR_3,
	h2f_ARLEN_0,
	nxt_in_ready,
	in_ready_hold,
	stateST_COMP_TRANS,
	out_valid_reg1,
	in_narrow_reg1,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	in_data_reg_68,
	cp_ready,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready1,
	sink0_data,
	Equal16,
	altera_reset_synchronizer_int_chain_out,
	in_data_reg_0,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	Add2,
	Add21,
	Add22,
	Add23,
	nxt_out_eop,
	Equal5,
	src1_valid,
	src_valid,
	cp_ready1,
	in_data_reg_69,
	src_valid1,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_6,
	sink0_endofpacket,
	write_cp_data_77,
	write_cp_data_78,
	write_cp_data_75,
	write_cp_data_74,
	write_cp_data_76,
	WideNor0,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	Selector3,
	Selector10,
	base_address_3,
	Selector4,
	Selector11,
	base_address_2,
	Selector5,
	Selector12,
	out_data_1,
	out_data_0,
	Selector6,
	Selector13,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARADDR_0;
input 	h2f_ARADDR_1;
input 	h2f_ARADDR_2;
input 	h2f_ARADDR_3;
input 	h2f_ARLEN_0;
output 	nxt_in_ready;
input 	in_ready_hold;
output 	stateST_COMP_TRANS;
output 	out_valid_reg1;
output 	in_narrow_reg1;
output 	in_byteen_reg_3;
output 	in_byteen_reg_2;
output 	in_byteen_reg_1;
output 	in_byteen_reg_0;
output 	in_data_reg_68;
input 	cp_ready;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready1;
input 	[128:0] sink0_data;
input 	Equal16;
input 	altera_reset_synchronizer_int_chain_out;
output 	in_data_reg_0;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
input 	Add2;
input 	Add21;
input 	Add22;
input 	Add23;
output 	nxt_out_eop;
input 	Equal5;
input 	src1_valid;
input 	src_valid;
input 	cp_ready1;
output 	in_data_reg_69;
input 	src_valid1;
output 	out_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_6;
input 	sink0_endofpacket;
input 	write_cp_data_77;
input 	write_cp_data_78;
input 	write_cp_data_75;
input 	write_cp_data_74;
input 	write_cp_data_76;
input 	WideNor0;
output 	in_data_reg_105;
output 	in_data_reg_106;
output 	in_data_reg_107;
output 	in_data_reg_108;
output 	in_data_reg_109;
output 	in_data_reg_110;
output 	in_data_reg_111;
output 	in_data_reg_112;
output 	in_data_reg_113;
output 	in_data_reg_114;
output 	in_data_reg_115;
output 	in_data_reg_116;
input 	Selector3;
input 	Selector10;
input 	base_address_3;
input 	Selector4;
input 	Selector11;
input 	base_address_2;
input 	Selector5;
input 	Selector12;
input 	out_data_1;
input 	out_data_0;
input 	Selector6;
input 	Selector13;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \align_address_to_size|LessThan0~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt[3]~1_combout ;
wire \nxt_uncomp_subburst_byte_cnt[4]~2_combout ;
wire \Add4~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt[5]~3_combout ;
wire \nxt_uncomp_subburst_byte_cnt[2]~4_combout ;
wire \nxt_uncomp_subburst_byte_cnt[6]~5_combout ;
wire \WideOr0~combout ;
wire \in_valid~combout ;
wire \Selector0~0_combout ;
wire \load_next_out_cmd~combout ;
wire \state.ST_IDLE~q ;
wire \Selector2~0_combout ;
wire \Selector2~1_combout ;
wire \Selector2~2_combout ;
wire \state.ST_UNCOMP_TRANS~q ;
wire \Selector1~2_combout ;
wire \Selector1~0_combout ;
wire \Selector1~3_combout ;
wire \int_bytes_remaining_reg[5]~q ;
wire \d0_int_bytes_remaining[2]~6_combout ;
wire \d0_int_bytes_remaining[2]~7_combout ;
wire \int_bytes_remaining_reg[2]~q ;
wire \d0_int_bytes_remaining[3]~4_combout ;
wire \d0_int_bytes_remaining[3]~5_combout ;
wire \int_bytes_remaining_reg[3]~q ;
wire \Add1~1_combout ;
wire \d0_int_bytes_remaining[4]~8_combout ;
wire \int_bytes_remaining_reg[4]~q ;
wire \Add1~0_combout ;
wire \d0_int_bytes_remaining[5]~0_combout ;
wire \d0_int_bytes_remaining[5]~1_combout ;
wire \int_bytes_remaining_reg[6]~q ;
wire \d0_int_bytes_remaining[6]~2_combout ;
wire \d0_int_bytes_remaining[6]~3_combout ;
wire \Equal0~0_combout ;
wire \new_burst_reg~0_combout ;
wire \new_burst_reg~q ;
wire \Selector1~1_combout ;
wire \WideNor0~0_combout ;
wire \NON_PIPELINED_INPUTS.load_next_cmd~combout ;
wire \in_bytecount_reg_zero~q ;
wire \nxt_out_valid~0_combout ;
wire \LessThan0~0_combout ;
wire \Selector3~0_combout ;
wire \in_size_reg[0]~q ;
wire \in_size_reg[2]~q ;
wire \in_size_reg[1]~q ;
wire \ShiftLeft0~0_combout ;
wire \ShiftLeft0~1_combout ;
wire \int_byte_cnt_narrow_reg[3]~q ;
wire \ShiftLeft0~2_combout ;
wire \int_byte_cnt_narrow_reg[2]~q ;
wire \ShiftLeft0~3_combout ;
wire \ShiftLeft0~4_combout ;
wire \int_byte_cnt_narrow_reg[1]~q ;
wire \int_byte_cnt_narrow_reg[0]~q ;
wire \Add0~13_sumout ;
wire \d0_int_nxt_addr[0]~3_combout ;
wire \in_burstwrap_reg[0]~q ;
wire \nxt_addr[0]~0_combout ;
wire \int_nxt_addr_reg[0]~q ;
wire \d0_int_nxt_addr[0]~4_combout ;
wire \int_nxt_addr_reg_dly[0]~q ;
wire \Add0~14 ;
wire \Add0~9_sumout ;
wire \in_burstwrap_reg[1]~q ;
wire \nxt_addr[1]~4_combout ;
wire \int_nxt_addr_reg[1]~q ;
wire \d0_int_nxt_addr[1]~7_combout ;
wire \d0_int_nxt_addr[1]~2_combout ;
wire \int_nxt_addr_reg_dly[1]~q ;
wire \Add0~10 ;
wire \Add0~6 ;
wire \Add0~1_sumout ;
wire \in_burstwrap_reg[3]~q ;
wire \nxt_addr[3]~12_combout ;
wire \int_nxt_addr_reg[3]~q ;
wire \d0_int_nxt_addr[3]~5_combout ;
wire \d0_int_nxt_addr[3]~0_combout ;
wire \Add0~5_sumout ;
wire \in_burstwrap_reg[2]~q ;
wire \nxt_addr[2]~8_combout ;
wire \int_nxt_addr_reg[2]~q ;
wire \d0_int_nxt_addr[2]~6_combout ;
wire \d0_int_nxt_addr[2]~1_combout ;
wire \in_eop_reg~q ;


spw_babasu_altera_merlin_address_alignment_6 align_address_to_size(
	.new_burst_reg(\new_burst_reg~q ),
	.src_data_86(sink0_data[86]),
	.in_size_reg_0(\in_size_reg[0]~q ),
	.ShiftLeft0(\ShiftLeft0~3_combout ),
	.LessThan0(\align_address_to_size|LessThan0~0_combout ));

cyclonev_lcell_comb \nxt_in_ready~1 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!in_ready_hold),
	.datac(!out_valid_reg1),
	.datad(!cp_ready),
	.datae(!stateST_COMP_TRANS),
	.dataf(!\new_burst_reg~q ),
	.datag(!stateST_UNCOMP_WR_SUBBURST),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~1 .extended_lut = "on";
defparam \nxt_in_ready~1 .lut_mask = 64'h2020F0F02020F0FF;
defparam \nxt_in_ready~1 .shared_arith = "off";

dffeas \state.ST_COMP_TRANS (
	.clk(clk_clk),
	.d(\Selector1~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_COMP_TRANS),
	.prn(vcc));
defparam \state.ST_COMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_COMP_TRANS .power_up = "low";

dffeas out_valid_reg(
	.clk(clk_clk),
	.d(\nxt_out_valid~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_valid_reg1),
	.prn(vcc));
defparam out_valid_reg.is_wysiwyg = "true";
defparam out_valid_reg.power_up = "low";

dffeas in_narrow_reg(
	.clk(clk_clk),
	.d(\LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_narrow_reg1),
	.prn(vcc));
defparam in_narrow_reg.is_wysiwyg = "true";
defparam in_narrow_reg.power_up = "low";

dffeas \in_byteen_reg[3] (
	.clk(clk_clk),
	.d(sink0_data[35]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_3),
	.prn(vcc));
defparam \in_byteen_reg[3] .is_wysiwyg = "true";
defparam \in_byteen_reg[3] .power_up = "low";

dffeas \in_byteen_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[34]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_2),
	.prn(vcc));
defparam \in_byteen_reg[2] .is_wysiwyg = "true";
defparam \in_byteen_reg[2] .power_up = "low";

dffeas \in_byteen_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[33]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_1),
	.prn(vcc));
defparam \in_byteen_reg[1] .is_wysiwyg = "true";
defparam \in_byteen_reg[1] .power_up = "low";

dffeas \in_byteen_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[32]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_0),
	.prn(vcc));
defparam \in_byteen_reg[0] .is_wysiwyg = "true";
defparam \in_byteen_reg[0] .power_up = "low";

dffeas \in_data_reg[68] (
	.clk(clk_clk),
	.d(sink0_data[68]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_68),
	.prn(vcc));
defparam \in_data_reg[68] .is_wysiwyg = "true";
defparam \in_data_reg[68] .power_up = "low";

dffeas \state.ST_UNCOMP_WR_SUBBURST (
	.clk(clk_clk),
	.d(\Selector3~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_UNCOMP_WR_SUBBURST),
	.prn(vcc));
defparam \state.ST_UNCOMP_WR_SUBBURST .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_WR_SUBBURST .power_up = "low";

cyclonev_lcell_comb \nxt_in_ready~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!out_valid_reg1),
	.datac(!cp_ready),
	.datad(!\state.ST_UNCOMP_TRANS~q ),
	.datae(!stateST_UNCOMP_WR_SUBBURST),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~0 .extended_lut = "off";
defparam \nxt_in_ready~0 .lut_mask = 64'h008A8A8A008A8A8A;
defparam \nxt_in_ready~0 .shared_arith = "off";

dffeas \in_data_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[0]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_0),
	.prn(vcc));
defparam \in_data_reg[0] .is_wysiwyg = "true";
defparam \in_data_reg[0] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[3] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[3]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_3),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[3] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[2] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[2]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_2),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[2] .power_up = "low";

cyclonev_lcell_comb \nxt_out_eop~0 (
	.dataa(!\in_eop_reg~q ),
	.datab(!stateST_COMP_TRANS),
	.datac(!\new_burst_reg~q ),
	.datad(!cp_ready),
	.datae(!\in_bytecount_reg_zero~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_out_eop),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_eop~0 .extended_lut = "off";
defparam \nxt_out_eop~0 .lut_mask = 64'h4447774744477747;
defparam \nxt_out_eop~0 .shared_arith = "off";

dffeas \in_data_reg[69] (
	.clk(clk_clk),
	.d(sink0_data[69]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_69),
	.prn(vcc));
defparam \in_data_reg[69] .is_wysiwyg = "true";
defparam \in_data_reg[69] .power_up = "low";

dffeas \out_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[3] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[3]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_3),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[3] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[3] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[2]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[4] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[4]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_4),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[4] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[4] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[5] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[5]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_5),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[5] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[5] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[6] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[6]~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_6),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[6] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[6] .power_up = "low";

dffeas \in_data_reg[105] (
	.clk(clk_clk),
	.d(sink0_data[105]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_105),
	.prn(vcc));
defparam \in_data_reg[105] .is_wysiwyg = "true";
defparam \in_data_reg[105] .power_up = "low";

dffeas \in_data_reg[106] (
	.clk(clk_clk),
	.d(sink0_data[106]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_106),
	.prn(vcc));
defparam \in_data_reg[106] .is_wysiwyg = "true";
defparam \in_data_reg[106] .power_up = "low";

dffeas \in_data_reg[107] (
	.clk(clk_clk),
	.d(sink0_data[107]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_107),
	.prn(vcc));
defparam \in_data_reg[107] .is_wysiwyg = "true";
defparam \in_data_reg[107] .power_up = "low";

dffeas \in_data_reg[108] (
	.clk(clk_clk),
	.d(sink0_data[108]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_108),
	.prn(vcc));
defparam \in_data_reg[108] .is_wysiwyg = "true";
defparam \in_data_reg[108] .power_up = "low";

dffeas \in_data_reg[109] (
	.clk(clk_clk),
	.d(sink0_data[109]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_109),
	.prn(vcc));
defparam \in_data_reg[109] .is_wysiwyg = "true";
defparam \in_data_reg[109] .power_up = "low";

dffeas \in_data_reg[110] (
	.clk(clk_clk),
	.d(sink0_data[110]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_110),
	.prn(vcc));
defparam \in_data_reg[110] .is_wysiwyg = "true";
defparam \in_data_reg[110] .power_up = "low";

dffeas \in_data_reg[111] (
	.clk(clk_clk),
	.d(sink0_data[111]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_111),
	.prn(vcc));
defparam \in_data_reg[111] .is_wysiwyg = "true";
defparam \in_data_reg[111] .power_up = "low";

dffeas \in_data_reg[112] (
	.clk(clk_clk),
	.d(sink0_data[112]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_112),
	.prn(vcc));
defparam \in_data_reg[112] .is_wysiwyg = "true";
defparam \in_data_reg[112] .power_up = "low";

dffeas \in_data_reg[113] (
	.clk(clk_clk),
	.d(sink0_data[113]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_113),
	.prn(vcc));
defparam \in_data_reg[113] .is_wysiwyg = "true";
defparam \in_data_reg[113] .power_up = "low";

dffeas \in_data_reg[114] (
	.clk(clk_clk),
	.d(sink0_data[114]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_114),
	.prn(vcc));
defparam \in_data_reg[114] .is_wysiwyg = "true";
defparam \in_data_reg[114] .power_up = "low";

dffeas \in_data_reg[115] (
	.clk(clk_clk),
	.d(sink0_data[115]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_115),
	.prn(vcc));
defparam \in_data_reg[115] .is_wysiwyg = "true";
defparam \in_data_reg[115] .power_up = "low";

dffeas \in_data_reg[116] (
	.clk(clk_clk),
	.d(sink0_data[116]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_116),
	.prn(vcc));
defparam \in_data_reg[116] .is_wysiwyg = "true";
defparam \in_data_reg[116] .power_up = "low";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt~0 (
	.dataa(!out_valid_reg1),
	.datab(!cp_ready),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt~0 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt~0 .lut_mask = 64'h1111111111111111;
defparam \nxt_uncomp_subburst_byte_cnt~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[3]~1 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!out_uncomp_byte_cnt_reg_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[3]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[3]~1 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[3]~1 .lut_mask = 64'h0FE40F4E0FE40F4E;
defparam \nxt_uncomp_subburst_byte_cnt[3]~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[4]~2 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!out_uncomp_byte_cnt_reg_2),
	.dataf(!out_uncomp_byte_cnt_reg_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[4]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[4]~2 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[4]~2 .lut_mask = 64'h00E40044FF4EFFEE;
defparam \nxt_uncomp_subburst_byte_cnt[4]~2 .shared_arith = "off";

cyclonev_lcell_comb \Add4~0 (
	.dataa(!out_uncomp_byte_cnt_reg_3),
	.datab(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datac(!out_uncomp_byte_cnt_reg_2),
	.datad(!out_uncomp_byte_cnt_reg_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add4~0 .extended_lut = "off";
defparam \Add4~0 .lut_mask = 64'h2000200020002000;
defparam \Add4~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[5]~3 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_5),
	.datae(!\Add4~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[5]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[5]~3 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[5]~3 .lut_mask = 64'h04FEAE5404FEAE54;
defparam \nxt_uncomp_subburst_byte_cnt[5]~3 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[2]~4 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[2]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[2]~4 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[2]~4 .lut_mask = 64'h0EF40EF40EF40EF4;
defparam \nxt_uncomp_subburst_byte_cnt[2]~4 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[6]~5 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_5),
	.datae(!\Add4~0_combout ),
	.dataf(!out_uncomp_byte_cnt_reg_6),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[6]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[6]~5 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[6]~5 .lut_mask = 64'h0404AE04FEFE54FE;
defparam \nxt_uncomp_subburst_byte_cnt[6]~5 .shared_arith = "off";

cyclonev_lcell_comb WideOr0(
	.dataa(!\nxt_uncomp_subburst_byte_cnt[3]~1_combout ),
	.datab(!\nxt_uncomp_subburst_byte_cnt[4]~2_combout ),
	.datac(!\nxt_uncomp_subburst_byte_cnt[5]~3_combout ),
	.datad(!\nxt_uncomp_subburst_byte_cnt[2]~4_combout ),
	.datae(!\nxt_uncomp_subburst_byte_cnt[6]~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr0.extended_lut = "off";
defparam WideOr0.lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam WideOr0.shared_arith = "off";

cyclonev_lcell_comb in_valid(
	.dataa(!in_ready_hold),
	.datab(!Equal16),
	.datac(!Equal5),
	.datad(!sink0_data[68]),
	.datae(!src1_valid),
	.dataf(!src_valid),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\in_valid~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam in_valid.extended_lut = "off";
defparam in_valid.lut_mask = 64'h0000000155555555;
defparam in_valid.shared_arith = "off";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!sink0_data[69]),
	.datab(!nxt_out_eop),
	.datac(!sink0_data[68]),
	.datad(!\in_valid~combout ),
	.datae(!\state.ST_IDLE~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'h005FCCFF005FCCFF;
defparam \Selector0~0 .shared_arith = "off";

cyclonev_lcell_comb load_next_out_cmd(
	.dataa(!out_valid_reg1),
	.datab(!cp_ready),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\load_next_out_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam load_next_out_cmd.extended_lut = "off";
defparam load_next_out_cmd.lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam load_next_out_cmd.shared_arith = "off";

dffeas \state.ST_IDLE (
	.clk(clk_clk),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_IDLE~q ),
	.prn(vcc));
defparam \state.ST_IDLE .is_wysiwyg = "true";
defparam \state.ST_IDLE .power_up = "low";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!nxt_out_eop),
	.datac(!stateST_UNCOMP_WR_SUBBURST),
	.datad(!\state.ST_IDLE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'h00EC00EC00EC00EC;
defparam \Selector2~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~1 (
	.dataa(!in_ready_hold),
	.datab(!Equal16),
	.datac(!Equal5),
	.datad(!sink0_data[68]),
	.datae(!src1_valid),
	.dataf(!\Selector2~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~1 .extended_lut = "off";
defparam \Selector2~1 .lut_mask = 64'h0000000100000000;
defparam \Selector2~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~2 (
	.dataa(!\WideOr0~combout ),
	.datab(!\Selector2~1_combout ),
	.datac(!\in_valid~combout ),
	.datad(!nxt_out_eop),
	.datae(!\state.ST_UNCOMP_TRANS~q ),
	.dataf(!sink0_data[69]),
	.datag(!stateST_UNCOMP_WR_SUBBURST),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~2 .extended_lut = "on";
defparam \Selector2~2 .lut_mask = 64'h3B33BB3F0A00AA00;
defparam \Selector2~2 .shared_arith = "off";

dffeas \state.ST_UNCOMP_TRANS (
	.clk(clk_clk),
	.d(\Selector2~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_UNCOMP_TRANS~q ),
	.prn(vcc));
defparam \state.ST_UNCOMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_TRANS .power_up = "low";

cyclonev_lcell_comb \Selector1~2 (
	.dataa(!in_ready_hold),
	.datab(!stateST_COMP_TRANS),
	.datac(!nxt_out_eop),
	.datad(!sink0_data[68]),
	.datae(gnd),
	.dataf(!src_valid),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~2 .extended_lut = "off";
defparam \Selector1~2 .lut_mask = 64'h3030303031303130;
defparam \Selector1~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!nxt_out_eop),
	.datac(!\state.ST_UNCOMP_TRANS~q ),
	.datad(!stateST_UNCOMP_WR_SUBBURST),
	.datae(!\state.ST_IDLE~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'h0000A8880000A888;
defparam \Selector1~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~3 (
	.dataa(!in_ready_hold),
	.datab(!sink0_data[69]),
	.datac(!src_valid),
	.datad(!src_valid1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~3 .extended_lut = "off";
defparam \Selector1~3 .lut_mask = 64'h0111011101110111;
defparam \Selector1~3 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[5] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[5]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[5]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[5] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[5] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[2]~6 (
	.dataa(!h2f_ARLEN_0),
	.datab(!sink0_data[69]),
	.datac(!sink0_data[68]),
	.datad(!write_cp_data_74),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[2]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[2]~6 .extended_lut = "off";
defparam \d0_int_bytes_remaining[2]~6 .lut_mask = 64'h2F222F222F222F22;
defparam \d0_int_bytes_remaining[2]~6 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[2]~7 (
	.dataa(!\new_burst_reg~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\int_bytes_remaining_reg[2]~q ),
	.datad(!\d0_int_bytes_remaining[2]~6_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[2]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[2]~7 .extended_lut = "off";
defparam \d0_int_bytes_remaining[2]~7 .lut_mask = 64'h287D287D287D287D;
defparam \d0_int_bytes_remaining[2]~7 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[2] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[2]~7_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[2]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[2] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[3]~4 (
	.dataa(!sink0_data[69]),
	.datab(!sink0_data[68]),
	.datac(!write_cp_data_75),
	.datad(!Add2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[3]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[3]~4 .extended_lut = "off";
defparam \d0_int_bytes_remaining[3]~4 .lut_mask = 64'h0357035703570357;
defparam \d0_int_bytes_remaining[3]~4 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[3]~5 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\int_bytes_remaining_reg[3]~q ),
	.datac(!out_byte_cnt_reg_2),
	.datad(!\int_bytes_remaining_reg[2]~q ),
	.datae(!\d0_int_bytes_remaining[3]~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[3]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[3]~5 .extended_lut = "off";
defparam \d0_int_bytes_remaining[3]~5 .lut_mask = 64'h28227D7728227D77;
defparam \d0_int_bytes_remaining[3]~5 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[3] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[3]~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[3]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[3] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[3] .power_up = "low";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!\int_bytes_remaining_reg[3]~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\int_bytes_remaining_reg[2]~q ),
	.datad(!\int_bytes_remaining_reg[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'hDF20DF20DF20DF20;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[4]~8 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!sink0_data[68]),
	.datad(!write_cp_data_76),
	.datae(!Add21),
	.dataf(!\Add1~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[4]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[4]~8 .extended_lut = "off";
defparam \d0_int_bytes_remaining[4]~8 .lut_mask = 64'hCCCFDDDF00031113;
defparam \d0_int_bytes_remaining[4]~8 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[4] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[4]~8_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[4]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[4] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[4] .power_up = "low";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!\int_bytes_remaining_reg[3]~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\int_bytes_remaining_reg[2]~q ),
	.datad(!\int_bytes_remaining_reg[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h2000200020002000;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[5]~0 (
	.dataa(!sink0_data[69]),
	.datab(!sink0_data[68]),
	.datac(!write_cp_data_77),
	.datad(!Add22),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[5]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[5]~0 .extended_lut = "off";
defparam \d0_int_bytes_remaining[5]~0 .lut_mask = 64'h0357035703570357;
defparam \d0_int_bytes_remaining[5]~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[5]~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\int_bytes_remaining_reg[5]~q ),
	.datac(!\Add1~0_combout ),
	.datad(!\d0_int_bytes_remaining[5]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[5]~1 .extended_lut = "off";
defparam \d0_int_bytes_remaining[5]~1 .lut_mask = 64'h287D287D287D287D;
defparam \d0_int_bytes_remaining[5]~1 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[6] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[6]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[6]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[6] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[6] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[6]~2 (
	.dataa(!sink0_data[69]),
	.datab(!sink0_data[68]),
	.datac(!write_cp_data_78),
	.datad(!Add23),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[6]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[6]~2 .extended_lut = "off";
defparam \d0_int_bytes_remaining[6]~2 .lut_mask = 64'h0357035703570357;
defparam \d0_int_bytes_remaining[6]~2 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[6]~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\int_bytes_remaining_reg[5]~q ),
	.datac(!\Add1~0_combout ),
	.datad(!\int_bytes_remaining_reg[6]~q ),
	.datae(!\d0_int_bytes_remaining[6]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[6]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[6]~3 .extended_lut = "off";
defparam \d0_int_bytes_remaining[6]~3 .lut_mask = 64'h08A25DF708A25DF7;
defparam \d0_int_bytes_remaining[6]~3 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!\d0_int_bytes_remaining[3]~5_combout ),
	.datab(!\d0_int_bytes_remaining[2]~7_combout ),
	.datac(!\d0_int_bytes_remaining[4]~8_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'h2020202020202020;
defparam \Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \new_burst_reg~0 (
	.dataa(!\Selector1~2_combout ),
	.datab(!\Selector1~0_combout ),
	.datac(!\Selector1~3_combout ),
	.datad(!\d0_int_bytes_remaining[5]~1_combout ),
	.datae(!\d0_int_bytes_remaining[6]~3_combout ),
	.dataf(!\Equal0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\new_burst_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \new_burst_reg~0 .extended_lut = "off";
defparam \new_burst_reg~0 .lut_mask = 64'hA2A2A2A2FFA2A2A2;
defparam \new_burst_reg~0 .shared_arith = "off";

dffeas new_burst_reg(
	.clk(clk_clk),
	.d(\new_burst_reg~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\new_burst_reg~q ),
	.prn(vcc));
defparam new_burst_reg.is_wysiwyg = "true";
defparam new_burst_reg.power_up = "low";

cyclonev_lcell_comb \Selector1~1 (
	.dataa(!sink0_data[69]),
	.datab(!stateST_COMP_TRANS),
	.datac(!nxt_out_eop),
	.datad(!sink0_data[68]),
	.datae(!\in_valid~combout ),
	.dataf(!\Selector1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~1 .extended_lut = "off";
defparam \Selector1~1 .lut_mask = 64'h3030777530303330;
defparam \Selector1~1 .shared_arith = "off";

cyclonev_lcell_comb \WideNor0~0 (
	.dataa(!sink0_data[69]),
	.datab(!sink0_data[68]),
	.datac(!WideNor0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideNor0~0 .extended_lut = "off";
defparam \WideNor0~0 .lut_mask = 64'h8A8A8A8A8A8A8A8A;
defparam \WideNor0~0 .shared_arith = "off";

cyclonev_lcell_comb \NON_PIPELINED_INPUTS.load_next_cmd (
	.dataa(!in_ready_hold),
	.datab(!nxt_in_ready1),
	.datac(!nxt_in_ready),
	.datad(!src_valid),
	.datae(!src_valid1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \NON_PIPELINED_INPUTS.load_next_cmd .extended_lut = "off";
defparam \NON_PIPELINED_INPUTS.load_next_cmd .lut_mask = 64'h0015151500151515;
defparam \NON_PIPELINED_INPUTS.load_next_cmd .shared_arith = "off";

dffeas in_bytecount_reg_zero(
	.clk(clk_clk),
	.d(\WideNor0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_bytecount_reg_zero~q ),
	.prn(vcc));
defparam in_bytecount_reg_zero.is_wysiwyg = "true";
defparam in_bytecount_reg_zero.power_up = "low";

cyclonev_lcell_comb \nxt_out_valid~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!\new_burst_reg~q ),
	.datac(!\in_bytecount_reg_zero~q ),
	.datad(!\in_valid~combout ),
	.datae(!cp_ready1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_valid~0 .extended_lut = "off";
defparam \nxt_out_valid~0 .lut_mask = 64'h50FF44FF50FF44FF;
defparam \nxt_out_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!sink0_data[87]),
	.datab(!sink0_data[88]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h8888888888888888;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~0 (
	.dataa(!nxt_out_eop),
	.datab(!\state.ST_UNCOMP_TRANS~q ),
	.datac(!stateST_UNCOMP_WR_SUBBURST),
	.datad(!\WideOr0~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'h002A002A002A002A;
defparam \Selector3~0 .shared_arith = "off";

dffeas \in_size_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[86]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[0]~q ),
	.prn(vcc));
defparam \in_size_reg[0] .is_wysiwyg = "true";
defparam \in_size_reg[0] .power_up = "low";

dffeas \in_size_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[88]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[2]~q ),
	.prn(vcc));
defparam \in_size_reg[2] .is_wysiwyg = "true";
defparam \in_size_reg[2] .power_up = "low";

dffeas \in_size_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[87]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[1]~q ),
	.prn(vcc));
defparam \in_size_reg[1] .is_wysiwyg = "true";
defparam \in_size_reg[1] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[87]),
	.datac(!sink0_data[88]),
	.datad(!\in_size_reg[2]~q ),
	.datae(!\in_size_reg[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~0 .extended_lut = "off";
defparam \ShiftLeft0~0 .lut_mask = 64'h1010BA101010BA10;
defparam \ShiftLeft0~0 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~1 .extended_lut = "off";
defparam \ShiftLeft0~1 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~1 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[3] (
	.clk(clk_clk),
	.d(\ShiftLeft0~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[3]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[3] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[3] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~2 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~2 .extended_lut = "off";
defparam \ShiftLeft0~2 .lut_mask = 64'h00E400E400E400E4;
defparam \ShiftLeft0~2 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[2] (
	.clk(clk_clk),
	.d(\ShiftLeft0~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[2]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[2] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[2] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[87]),
	.datac(!sink0_data[88]),
	.datad(!\in_size_reg[2]~q ),
	.datae(!\in_size_reg[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~3 .extended_lut = "off";
defparam \ShiftLeft0~3 .lut_mask = 64'hEA404040EA404040;
defparam \ShiftLeft0~3 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~4 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~4 .extended_lut = "off";
defparam \ShiftLeft0~4 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~4 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[1] (
	.clk(clk_clk),
	.d(\ShiftLeft0~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[1]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[1] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[1] .power_up = "low";

dffeas \int_byte_cnt_narrow_reg[0] (
	.clk(clk_clk),
	.d(\align_address_to_size|LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[0]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[0] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[0] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[0]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~3 (
	.dataa(!h2f_ARADDR_0),
	.datab(!sink0_data[69]),
	.datac(!sink0_data[68]),
	.datad(!out_data_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~3 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~3 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[0]~3 .shared_arith = "off";

dffeas \in_burstwrap_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[79]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[0]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[0] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[0] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[0]~0 (
	.dataa(!Selector13),
	.datab(!Selector6),
	.datac(!sink0_data[68]),
	.datad(!sink0_data[69]),
	.datae(!\new_burst_reg~q ),
	.dataf(!\d0_int_nxt_addr[0]~4_combout ),
	.datag(!\in_burstwrap_reg[0]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[0]~0 .extended_lut = "on";
defparam \nxt_addr[0]~0 .lut_mask = 64'h00000000F0F0FCA8;
defparam \nxt_addr[0]~0 .shared_arith = "off";

dffeas \int_nxt_addr_reg[0] (
	.clk(clk_clk),
	.d(\nxt_addr[0]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[0] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~4 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\Add0~13_sumout ),
	.datac(!\align_address_to_size|LessThan0~0_combout ),
	.datad(!\d0_int_nxt_addr[0]~3_combout ),
	.datae(!\int_nxt_addr_reg[0]~q ),
	.dataf(!\in_burstwrap_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~4 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~4 .lut_mask = 64'h0005AAAF2227AAAF;
defparam \d0_int_nxt_addr[0]~4 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[0] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[0]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[0] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[1]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[1]~q ),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \in_burstwrap_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[80]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[1]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[1] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[1] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[1]~4 (
	.dataa(!Selector12),
	.datab(!Selector5),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!\new_burst_reg~q ),
	.dataf(!\d0_int_nxt_addr[1]~2_combout ),
	.datag(!\in_burstwrap_reg[1]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[1]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[1]~4 .extended_lut = "on";
defparam \nxt_addr[1]~4 .lut_mask = 64'h00000000F0F0FAC8;
defparam \nxt_addr[1]~4 .shared_arith = "off";

dffeas \int_nxt_addr_reg[1] (
	.clk(clk_clk),
	.d(\nxt_addr[1]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[1] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~7 (
	.dataa(!h2f_ARADDR_1),
	.datab(!sink0_data[69]),
	.datac(!sink0_data[68]),
	.datad(!out_data_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~7 .extended_lut = "off";
defparam \d0_int_nxt_addr[1]~7 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[1]~7 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~2 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\Add0~9_sumout ),
	.datac(!\in_burstwrap_reg[1]~q ),
	.datad(!\int_nxt_addr_reg[1]~q ),
	.datae(!\ShiftLeft0~3_combout ),
	.dataf(!\d0_int_nxt_addr[1]~7_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~2 .extended_lut = "off";
defparam \d0_int_nxt_addr[1]~2 .lut_mask = 64'h02AA02AA02AA57FF;
defparam \d0_int_nxt_addr[1]~2 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[1] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[1]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[1] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_2),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[2]~q ),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[3]~q ),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

dffeas \in_burstwrap_reg[3] (
	.clk(clk_clk),
	.d(sink0_data[82]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[3]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[3] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[3] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[3]~12 (
	.dataa(!Selector10),
	.datab(!Selector3),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!\new_burst_reg~q ),
	.dataf(!\d0_int_nxt_addr[3]~0_combout ),
	.datag(!\in_burstwrap_reg[3]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[3]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[3]~12 .extended_lut = "on";
defparam \nxt_addr[3]~12 .lut_mask = 64'h00000000F0F0FAC8;
defparam \nxt_addr[3]~12 .shared_arith = "off";

dffeas \int_nxt_addr_reg[3] (
	.clk(clk_clk),
	.d(\nxt_addr[3]~12_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[3]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[3] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~5 (
	.dataa(!\Add0~1_sumout ),
	.datab(!\in_burstwrap_reg[3]~q ),
	.datac(!\int_nxt_addr_reg[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~5 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~5 .lut_mask = 64'hE0E0E0E0E0E0E0E0;
defparam \d0_int_nxt_addr[3]~5 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!h2f_ARADDR_3),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!base_address_3),
	.dataf(!\d0_int_nxt_addr[3]~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~0 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~0 .lut_mask = 64'hABABABFF01010155;
defparam \d0_int_nxt_addr[3]~0 .shared_arith = "off";

dffeas \in_burstwrap_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[81]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[2]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[2] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[2] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[2]~8 (
	.dataa(!Selector11),
	.datab(!Selector4),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!\new_burst_reg~q ),
	.dataf(!\d0_int_nxt_addr[2]~1_combout ),
	.datag(!\in_burstwrap_reg[2]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[2]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[2]~8 .extended_lut = "on";
defparam \nxt_addr[2]~8 .lut_mask = 64'h00000000F0F0FAC8;
defparam \nxt_addr[2]~8 .shared_arith = "off";

dffeas \int_nxt_addr_reg[2] (
	.clk(clk_clk),
	.d(\nxt_addr[2]~8_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[2]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~6 (
	.dataa(!\Add0~5_sumout ),
	.datab(!\in_burstwrap_reg[2]~q ),
	.datac(!\int_nxt_addr_reg[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~6 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~6 .lut_mask = 64'hE0E0E0E0E0E0E0E0;
defparam \d0_int_nxt_addr[2]~6 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!h2f_ARADDR_2),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!base_address_2),
	.dataf(!\d0_int_nxt_addr[2]~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~1 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~1 .lut_mask = 64'hABABABFF01010155;
defparam \d0_int_nxt_addr[2]~1 .shared_arith = "off";

dffeas in_eop_reg(
	.clk(clk_clk),
	.d(sink0_endofpacket),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_eop_reg~q ),
	.prn(vcc));
defparam in_eop_reg.is_wysiwyg = "true";
defparam in_eop_reg.power_up = "low";

endmodule

module spw_babasu_altera_merlin_address_alignment_6 (
	new_burst_reg,
	src_data_86,
	in_size_reg_0,
	ShiftLeft0,
	LessThan0)/* synthesis synthesis_greybox=0 */;
input 	new_burst_reg;
input 	src_data_86;
input 	in_size_reg_0;
input 	ShiftLeft0;
output 	LessThan0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!new_burst_reg),
	.datab(!src_data_86),
	.datac(!in_size_reg_0),
	.datad(!ShiftLeft0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan0),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h00E400E400E400E4;
defparam \LessThan0~0 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_burst_adapter_6 (
	h2f_ARADDR_0,
	h2f_ARADDR_1,
	h2f_ARADDR_2,
	h2f_ARADDR_3,
	h2f_ARLEN_0,
	nxt_in_ready,
	in_ready_hold,
	saved_grant_1,
	stateST_COMP_TRANS,
	out_valid_reg,
	mem_used_1,
	in_narrow_reg,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	in_data_reg_68,
	cp_ready,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready1,
	sop_enable,
	saved_grant_0,
	altera_reset_synchronizer_int_chain_out,
	in_data_reg_0,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	Add2,
	Add21,
	Add22,
	Add23,
	burst_bytecount_5,
	write_cp_data_77,
	burst_bytecount_6,
	write_cp_data_78,
	burst_bytecount_3,
	write_cp_data_75,
	burst_bytecount_2,
	write_cp_data_74,
	burst_bytecount_4,
	write_cp_data_76,
	WideNor0,
	src0_valid,
	src0_valid1,
	nxt_in_ready2,
	src_valid,
	src_payload_0,
	nxt_out_eop,
	cp_ready1,
	in_data_reg_69,
	src_data_87,
	src_data_88,
	src_data_35,
	src_data_34,
	src_data_33,
	src_data_32,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_6,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	Selector3,
	Selector10,
	base_address_3,
	Selector4,
	Selector11,
	base_address_2,
	src_payload,
	src_data_82,
	src_data_81,
	src_data_105,
	src_data_106,
	src_data_107,
	src_data_108,
	src_data_109,
	src_data_110,
	src_data_111,
	src_data_112,
	src_data_113,
	src_data_114,
	src_data_115,
	src_data_116,
	src_data_86,
	Selector5,
	Selector12,
	out_data_1,
	src_data_80,
	out_data_0,
	Selector6,
	Selector13,
	src_data_79,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARADDR_0;
input 	h2f_ARADDR_1;
input 	h2f_ARADDR_2;
input 	h2f_ARADDR_3;
input 	h2f_ARLEN_0;
output 	nxt_in_ready;
input 	in_ready_hold;
input 	saved_grant_1;
output 	stateST_COMP_TRANS;
output 	out_valid_reg;
input 	mem_used_1;
output 	in_narrow_reg;
output 	in_byteen_reg_3;
output 	in_byteen_reg_2;
output 	in_byteen_reg_1;
output 	in_byteen_reg_0;
output 	in_data_reg_68;
input 	cp_ready;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready1;
input 	sop_enable;
input 	saved_grant_0;
input 	altera_reset_synchronizer_int_chain_out;
output 	in_data_reg_0;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
input 	Add2;
input 	Add21;
input 	Add22;
input 	Add23;
input 	burst_bytecount_5;
input 	write_cp_data_77;
input 	burst_bytecount_6;
input 	write_cp_data_78;
input 	burst_bytecount_3;
input 	write_cp_data_75;
input 	burst_bytecount_2;
input 	write_cp_data_74;
input 	burst_bytecount_4;
input 	write_cp_data_76;
output 	WideNor0;
input 	src0_valid;
input 	src0_valid1;
output 	nxt_in_ready2;
input 	src_valid;
input 	src_payload_0;
output 	nxt_out_eop;
input 	cp_ready1;
output 	in_data_reg_69;
input 	src_data_87;
input 	src_data_88;
input 	src_data_35;
input 	src_data_34;
input 	src_data_33;
input 	src_data_32;
output 	out_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_6;
output 	in_data_reg_105;
output 	in_data_reg_106;
output 	in_data_reg_107;
output 	in_data_reg_108;
output 	in_data_reg_109;
output 	in_data_reg_110;
output 	in_data_reg_111;
output 	in_data_reg_112;
output 	in_data_reg_113;
output 	in_data_reg_114;
output 	in_data_reg_115;
output 	in_data_reg_116;
input 	Selector3;
input 	Selector10;
input 	base_address_3;
input 	Selector4;
input 	Selector11;
input 	base_address_2;
input 	src_payload;
input 	src_data_82;
input 	src_data_81;
input 	src_data_105;
input 	src_data_106;
input 	src_data_107;
input 	src_data_108;
input 	src_data_109;
input 	src_data_110;
input 	src_data_111;
input 	src_data_112;
input 	src_data_113;
input 	src_data_114;
input 	src_data_115;
input 	src_data_116;
input 	src_data_86;
input 	Selector5;
input 	Selector12;
input 	out_data_1;
input 	src_data_80;
input 	out_data_0;
input 	Selector6;
input 	Selector13;
input 	src_data_79;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



spw_babasu_altera_merlin_burst_adapter_13_1_6 \altera_merlin_burst_adapter_13_1.burst_adapter (
	.h2f_ARADDR_0(h2f_ARADDR_0),
	.h2f_ARADDR_1(h2f_ARADDR_1),
	.h2f_ARADDR_2(h2f_ARADDR_2),
	.h2f_ARADDR_3(h2f_ARADDR_3),
	.h2f_ARLEN_0(h2f_ARLEN_0),
	.nxt_in_ready(nxt_in_ready),
	.in_ready_hold(in_ready_hold),
	.sink0_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_116,src_data_115,src_data_114,src_data_113,src_data_112,src_data_111,src_data_110,src_data_109,src_data_108,src_data_107,src_data_106,src_data_105,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_88,src_data_87,
src_data_86,gnd,gnd,gnd,src_data_82,src_data_81,src_data_80,src_data_79,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,saved_grant_1,saved_grant_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_35,src_data_34,src_data_33,
src_data_32,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_payload}),
	.stateST_COMP_TRANS(stateST_COMP_TRANS),
	.out_valid_reg1(out_valid_reg),
	.mem_used_1(mem_used_1),
	.in_narrow_reg1(in_narrow_reg),
	.in_byteen_reg_3(in_byteen_reg_3),
	.in_byteen_reg_2(in_byteen_reg_2),
	.in_byteen_reg_1(in_byteen_reg_1),
	.in_byteen_reg_0(in_byteen_reg_0),
	.in_data_reg_68(in_data_reg_68),
	.cp_ready(cp_ready),
	.stateST_UNCOMP_WR_SUBBURST(stateST_UNCOMP_WR_SUBBURST),
	.nxt_in_ready1(nxt_in_ready1),
	.sop_enable(sop_enable),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.in_data_reg_0(in_data_reg_0),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_3),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_2),
	.Add2(Add2),
	.Add21(Add21),
	.Add22(Add22),
	.Add23(Add23),
	.burst_bytecount_5(burst_bytecount_5),
	.write_cp_data_77(write_cp_data_77),
	.burst_bytecount_6(burst_bytecount_6),
	.write_cp_data_78(write_cp_data_78),
	.burst_bytecount_3(burst_bytecount_3),
	.write_cp_data_75(write_cp_data_75),
	.burst_bytecount_2(burst_bytecount_2),
	.write_cp_data_74(write_cp_data_74),
	.burst_bytecount_4(burst_bytecount_4),
	.write_cp_data_76(write_cp_data_76),
	.WideNor0(WideNor0),
	.src0_valid(src0_valid),
	.src0_valid1(src0_valid1),
	.nxt_in_ready2(nxt_in_ready2),
	.src_valid(src_valid),
	.sink0_endofpacket(src_payload_0),
	.nxt_out_eop(nxt_out_eop),
	.cp_ready1(cp_ready1),
	.in_data_reg_69(in_data_reg_69),
	.out_byte_cnt_reg_2(out_byte_cnt_reg_2),
	.out_uncomp_byte_cnt_reg_3(out_uncomp_byte_cnt_reg_3),
	.out_uncomp_byte_cnt_reg_2(out_uncomp_byte_cnt_reg_2),
	.out_uncomp_byte_cnt_reg_4(out_uncomp_byte_cnt_reg_4),
	.out_uncomp_byte_cnt_reg_5(out_uncomp_byte_cnt_reg_5),
	.out_uncomp_byte_cnt_reg_6(out_uncomp_byte_cnt_reg_6),
	.in_data_reg_105(in_data_reg_105),
	.in_data_reg_106(in_data_reg_106),
	.in_data_reg_107(in_data_reg_107),
	.in_data_reg_108(in_data_reg_108),
	.in_data_reg_109(in_data_reg_109),
	.in_data_reg_110(in_data_reg_110),
	.in_data_reg_111(in_data_reg_111),
	.in_data_reg_112(in_data_reg_112),
	.in_data_reg_113(in_data_reg_113),
	.in_data_reg_114(in_data_reg_114),
	.in_data_reg_115(in_data_reg_115),
	.in_data_reg_116(in_data_reg_116),
	.Selector3(Selector3),
	.Selector10(Selector10),
	.base_address_3(base_address_3),
	.Selector4(Selector4),
	.Selector11(Selector11),
	.base_address_2(base_address_2),
	.Selector5(Selector5),
	.Selector12(Selector12),
	.out_data_1(out_data_1),
	.out_data_0(out_data_0),
	.Selector6(Selector6),
	.Selector13(Selector13),
	.clk_clk(clk_clk));

endmodule

module spw_babasu_altera_merlin_burst_adapter_13_1_6 (
	h2f_ARADDR_0,
	h2f_ARADDR_1,
	h2f_ARADDR_2,
	h2f_ARADDR_3,
	h2f_ARLEN_0,
	nxt_in_ready,
	in_ready_hold,
	sink0_data,
	stateST_COMP_TRANS,
	out_valid_reg1,
	mem_used_1,
	in_narrow_reg1,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	in_data_reg_68,
	cp_ready,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready1,
	sop_enable,
	altera_reset_synchronizer_int_chain_out,
	in_data_reg_0,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	Add2,
	Add21,
	Add22,
	Add23,
	burst_bytecount_5,
	write_cp_data_77,
	burst_bytecount_6,
	write_cp_data_78,
	burst_bytecount_3,
	write_cp_data_75,
	burst_bytecount_2,
	write_cp_data_74,
	burst_bytecount_4,
	write_cp_data_76,
	WideNor0,
	src0_valid,
	src0_valid1,
	nxt_in_ready2,
	src_valid,
	sink0_endofpacket,
	nxt_out_eop,
	cp_ready1,
	in_data_reg_69,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_6,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	Selector3,
	Selector10,
	base_address_3,
	Selector4,
	Selector11,
	base_address_2,
	Selector5,
	Selector12,
	out_data_1,
	out_data_0,
	Selector6,
	Selector13,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARADDR_0;
input 	h2f_ARADDR_1;
input 	h2f_ARADDR_2;
input 	h2f_ARADDR_3;
input 	h2f_ARLEN_0;
output 	nxt_in_ready;
input 	in_ready_hold;
input 	[128:0] sink0_data;
output 	stateST_COMP_TRANS;
output 	out_valid_reg1;
input 	mem_used_1;
output 	in_narrow_reg1;
output 	in_byteen_reg_3;
output 	in_byteen_reg_2;
output 	in_byteen_reg_1;
output 	in_byteen_reg_0;
output 	in_data_reg_68;
input 	cp_ready;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready1;
input 	sop_enable;
input 	altera_reset_synchronizer_int_chain_out;
output 	in_data_reg_0;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
input 	Add2;
input 	Add21;
input 	Add22;
input 	Add23;
input 	burst_bytecount_5;
input 	write_cp_data_77;
input 	burst_bytecount_6;
input 	write_cp_data_78;
input 	burst_bytecount_3;
input 	write_cp_data_75;
input 	burst_bytecount_2;
input 	write_cp_data_74;
input 	burst_bytecount_4;
input 	write_cp_data_76;
output 	WideNor0;
input 	src0_valid;
input 	src0_valid1;
output 	nxt_in_ready2;
input 	src_valid;
input 	sink0_endofpacket;
output 	nxt_out_eop;
input 	cp_ready1;
output 	in_data_reg_69;
output 	out_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_6;
output 	in_data_reg_105;
output 	in_data_reg_106;
output 	in_data_reg_107;
output 	in_data_reg_108;
output 	in_data_reg_109;
output 	in_data_reg_110;
output 	in_data_reg_111;
output 	in_data_reg_112;
output 	in_data_reg_113;
output 	in_data_reg_114;
output 	in_data_reg_115;
output 	in_data_reg_116;
input 	Selector3;
input 	Selector10;
input 	base_address_3;
input 	Selector4;
input 	Selector11;
input 	base_address_2;
input 	Selector5;
input 	Selector12;
input 	out_data_1;
input 	out_data_0;
input 	Selector6;
input 	Selector13;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \align_address_to_size|LessThan0~0_combout ;
wire \nxt_in_ready~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt[3]~1_combout ;
wire \nxt_uncomp_subburst_byte_cnt[4]~2_combout ;
wire \Add4~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt[5]~3_combout ;
wire \nxt_uncomp_subburst_byte_cnt[2]~4_combout ;
wire \nxt_uncomp_subburst_byte_cnt[6]~5_combout ;
wire \WideOr0~combout ;
wire \Selector2~0_combout ;
wire \nxt_in_ready~3_combout ;
wire \Selector0~0_combout ;
wire \Selector0~1_combout ;
wire \Selector0~2_combout ;
wire \load_next_out_cmd~combout ;
wire \state.ST_IDLE~q ;
wire \Selector2~1_combout ;
wire \Selector2~2_combout ;
wire \state.ST_UNCOMP_TRANS~q ;
wire \in_valid~combout ;
wire \Selector1~0_combout ;
wire \Selector1~1_combout ;
wire \int_bytes_remaining_reg[5]~q ;
wire \d0_int_bytes_remaining[2]~4_combout ;
wire \d0_int_bytes_remaining[2]~5_combout ;
wire \int_bytes_remaining_reg[2]~q ;
wire \d0_int_bytes_remaining[3]~6_combout ;
wire \d0_int_bytes_remaining[3]~7_combout ;
wire \int_bytes_remaining_reg[3]~q ;
wire \Add1~1_combout ;
wire \d0_int_bytes_remaining[4]~8_combout ;
wire \int_bytes_remaining_reg[4]~q ;
wire \Add1~0_combout ;
wire \d0_int_bytes_remaining[5]~0_combout ;
wire \d0_int_bytes_remaining[5]~1_combout ;
wire \int_bytes_remaining_reg[6]~q ;
wire \d0_int_bytes_remaining[6]~2_combout ;
wire \d0_int_bytes_remaining[6]~3_combout ;
wire \Equal0~0_combout ;
wire \new_burst_reg~0_combout ;
wire \new_burst_reg~q ;
wire \Selector1~2_combout ;
wire \WideNor0~1_combout ;
wire \NON_PIPELINED_INPUTS.load_next_cmd~combout ;
wire \in_bytecount_reg_zero~q ;
wire \nxt_out_valid~0_combout ;
wire \nxt_out_valid~1_combout ;
wire \LessThan0~0_combout ;
wire \Selector3~0_combout ;
wire \in_size_reg[0]~q ;
wire \in_size_reg[1]~q ;
wire \in_size_reg[2]~q ;
wire \ShiftLeft0~0_combout ;
wire \ShiftLeft0~1_combout ;
wire \int_byte_cnt_narrow_reg[3]~q ;
wire \ShiftLeft0~2_combout ;
wire \int_byte_cnt_narrow_reg[2]~q ;
wire \ShiftLeft0~3_combout ;
wire \ShiftLeft0~4_combout ;
wire \int_byte_cnt_narrow_reg[1]~q ;
wire \int_byte_cnt_narrow_reg[0]~q ;
wire \Add0~13_sumout ;
wire \d0_int_nxt_addr[0]~3_combout ;
wire \in_burstwrap_reg[0]~q ;
wire \nxt_addr[0]~0_combout ;
wire \int_nxt_addr_reg[0]~q ;
wire \d0_int_nxt_addr[0]~4_combout ;
wire \int_nxt_addr_reg_dly[0]~q ;
wire \Add0~14 ;
wire \Add0~9_sumout ;
wire \in_burstwrap_reg[1]~q ;
wire \nxt_addr[1]~4_combout ;
wire \int_nxt_addr_reg[1]~q ;
wire \d0_int_nxt_addr[1]~7_combout ;
wire \d0_int_nxt_addr[1]~2_combout ;
wire \int_nxt_addr_reg_dly[1]~q ;
wire \Add0~10 ;
wire \Add0~6 ;
wire \Add0~1_sumout ;
wire \in_burstwrap_reg[3]~q ;
wire \nxt_addr[3]~12_combout ;
wire \int_nxt_addr_reg[3]~q ;
wire \d0_int_nxt_addr[3]~5_combout ;
wire \d0_int_nxt_addr[3]~0_combout ;
wire \Add0~5_sumout ;
wire \in_burstwrap_reg[2]~q ;
wire \nxt_addr[2]~8_combout ;
wire \int_nxt_addr_reg[2]~q ;
wire \d0_int_nxt_addr[2]~6_combout ;
wire \d0_int_nxt_addr[2]~1_combout ;
wire \in_eop_reg~q ;


spw_babasu_altera_merlin_address_alignment_7 align_address_to_size(
	.new_burst_reg(\new_burst_reg~q ),
	.src_data_86(sink0_data[86]),
	.in_size_reg_0(\in_size_reg[0]~q ),
	.ShiftLeft0(\ShiftLeft0~3_combout ),
	.LessThan0(\align_address_to_size|LessThan0~0_combout ));

cyclonev_lcell_comb \nxt_in_ready~4 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!in_ready_hold),
	.datac(!out_valid_reg1),
	.datad(!cp_ready),
	.datae(!stateST_COMP_TRANS),
	.dataf(!\new_burst_reg~q ),
	.datag(!stateST_UNCOMP_WR_SUBBURST),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~4 .extended_lut = "on";
defparam \nxt_in_ready~4 .lut_mask = 64'h2020F0F02020F0FF;
defparam \nxt_in_ready~4 .shared_arith = "off";

dffeas \state.ST_COMP_TRANS (
	.clk(clk_clk),
	.d(\Selector1~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_COMP_TRANS),
	.prn(vcc));
defparam \state.ST_COMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_COMP_TRANS .power_up = "low";

dffeas out_valid_reg(
	.clk(clk_clk),
	.d(\nxt_out_valid~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_valid_reg1),
	.prn(vcc));
defparam out_valid_reg.is_wysiwyg = "true";
defparam out_valid_reg.power_up = "low";

dffeas in_narrow_reg(
	.clk(clk_clk),
	.d(\LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_narrow_reg1),
	.prn(vcc));
defparam in_narrow_reg.is_wysiwyg = "true";
defparam in_narrow_reg.power_up = "low";

dffeas \in_byteen_reg[3] (
	.clk(clk_clk),
	.d(sink0_data[35]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_3),
	.prn(vcc));
defparam \in_byteen_reg[3] .is_wysiwyg = "true";
defparam \in_byteen_reg[3] .power_up = "low";

dffeas \in_byteen_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[34]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_2),
	.prn(vcc));
defparam \in_byteen_reg[2] .is_wysiwyg = "true";
defparam \in_byteen_reg[2] .power_up = "low";

dffeas \in_byteen_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[33]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_1),
	.prn(vcc));
defparam \in_byteen_reg[1] .is_wysiwyg = "true";
defparam \in_byteen_reg[1] .power_up = "low";

dffeas \in_byteen_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[32]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_0),
	.prn(vcc));
defparam \in_byteen_reg[0] .is_wysiwyg = "true";
defparam \in_byteen_reg[0] .power_up = "low";

dffeas \in_data_reg[68] (
	.clk(clk_clk),
	.d(sink0_data[68]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_68),
	.prn(vcc));
defparam \in_data_reg[68] .is_wysiwyg = "true";
defparam \in_data_reg[68] .power_up = "low";

dffeas \state.ST_UNCOMP_WR_SUBBURST (
	.clk(clk_clk),
	.d(\Selector3~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_UNCOMP_WR_SUBBURST),
	.prn(vcc));
defparam \state.ST_UNCOMP_WR_SUBBURST .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_WR_SUBBURST .power_up = "low";

cyclonev_lcell_comb \nxt_in_ready~1 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!out_valid_reg1),
	.datac(!cp_ready),
	.datad(!\nxt_in_ready~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~1 .extended_lut = "off";
defparam \nxt_in_ready~1 .lut_mask = 64'h8A008A008A008A00;
defparam \nxt_in_ready~1 .shared_arith = "off";

dffeas \in_data_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[0]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_0),
	.prn(vcc));
defparam \in_data_reg[0] .is_wysiwyg = "true";
defparam \in_data_reg[0] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[3] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[3]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_3),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[3] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[2] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[2]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_2),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[2] .power_up = "low";

cyclonev_lcell_comb \WideNor0~0 (
	.dataa(!sop_enable),
	.datab(!burst_bytecount_2),
	.datac(!burst_bytecount_3),
	.datad(!burst_bytecount_4),
	.datae(!burst_bytecount_5),
	.dataf(!burst_bytecount_6),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideNor0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideNor0~0 .extended_lut = "off";
defparam \WideNor0~0 .lut_mask = 64'h4000000000000000;
defparam \WideNor0~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_in_ready~2 (
	.dataa(!nxt_in_ready1),
	.datab(!nxt_in_ready),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready2),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~2 .extended_lut = "off";
defparam \nxt_in_ready~2 .lut_mask = 64'h8888888888888888;
defparam \nxt_in_ready~2 .shared_arith = "off";

cyclonev_lcell_comb \nxt_out_eop~0 (
	.dataa(!\in_eop_reg~q ),
	.datab(!stateST_COMP_TRANS),
	.datac(!\new_burst_reg~q ),
	.datad(!cp_ready),
	.datae(!\in_bytecount_reg_zero~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_out_eop),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_eop~0 .extended_lut = "off";
defparam \nxt_out_eop~0 .lut_mask = 64'h4447774744477747;
defparam \nxt_out_eop~0 .shared_arith = "off";

dffeas \in_data_reg[69] (
	.clk(clk_clk),
	.d(sink0_data[69]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_69),
	.prn(vcc));
defparam \in_data_reg[69] .is_wysiwyg = "true";
defparam \in_data_reg[69] .power_up = "low";

dffeas \out_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[3] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[3]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_3),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[3] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[3] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[2]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[4] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[4]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_4),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[4] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[4] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[5] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[5]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_5),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[5] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[5] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[6] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[6]~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_6),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[6] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[6] .power_up = "low";

dffeas \in_data_reg[105] (
	.clk(clk_clk),
	.d(sink0_data[105]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_105),
	.prn(vcc));
defparam \in_data_reg[105] .is_wysiwyg = "true";
defparam \in_data_reg[105] .power_up = "low";

dffeas \in_data_reg[106] (
	.clk(clk_clk),
	.d(sink0_data[106]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_106),
	.prn(vcc));
defparam \in_data_reg[106] .is_wysiwyg = "true";
defparam \in_data_reg[106] .power_up = "low";

dffeas \in_data_reg[107] (
	.clk(clk_clk),
	.d(sink0_data[107]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_107),
	.prn(vcc));
defparam \in_data_reg[107] .is_wysiwyg = "true";
defparam \in_data_reg[107] .power_up = "low";

dffeas \in_data_reg[108] (
	.clk(clk_clk),
	.d(sink0_data[108]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_108),
	.prn(vcc));
defparam \in_data_reg[108] .is_wysiwyg = "true";
defparam \in_data_reg[108] .power_up = "low";

dffeas \in_data_reg[109] (
	.clk(clk_clk),
	.d(sink0_data[109]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_109),
	.prn(vcc));
defparam \in_data_reg[109] .is_wysiwyg = "true";
defparam \in_data_reg[109] .power_up = "low";

dffeas \in_data_reg[110] (
	.clk(clk_clk),
	.d(sink0_data[110]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_110),
	.prn(vcc));
defparam \in_data_reg[110] .is_wysiwyg = "true";
defparam \in_data_reg[110] .power_up = "low";

dffeas \in_data_reg[111] (
	.clk(clk_clk),
	.d(sink0_data[111]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_111),
	.prn(vcc));
defparam \in_data_reg[111] .is_wysiwyg = "true";
defparam \in_data_reg[111] .power_up = "low";

dffeas \in_data_reg[112] (
	.clk(clk_clk),
	.d(sink0_data[112]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_112),
	.prn(vcc));
defparam \in_data_reg[112] .is_wysiwyg = "true";
defparam \in_data_reg[112] .power_up = "low";

dffeas \in_data_reg[113] (
	.clk(clk_clk),
	.d(sink0_data[113]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_113),
	.prn(vcc));
defparam \in_data_reg[113] .is_wysiwyg = "true";
defparam \in_data_reg[113] .power_up = "low";

dffeas \in_data_reg[114] (
	.clk(clk_clk),
	.d(sink0_data[114]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_114),
	.prn(vcc));
defparam \in_data_reg[114] .is_wysiwyg = "true";
defparam \in_data_reg[114] .power_up = "low";

dffeas \in_data_reg[115] (
	.clk(clk_clk),
	.d(sink0_data[115]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_115),
	.prn(vcc));
defparam \in_data_reg[115] .is_wysiwyg = "true";
defparam \in_data_reg[115] .power_up = "low";

dffeas \in_data_reg[116] (
	.clk(clk_clk),
	.d(sink0_data[116]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_116),
	.prn(vcc));
defparam \in_data_reg[116] .is_wysiwyg = "true";
defparam \in_data_reg[116] .power_up = "low";

cyclonev_lcell_comb \nxt_in_ready~0 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_in_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~0 .extended_lut = "off";
defparam \nxt_in_ready~0 .lut_mask = 64'h8888888888888888;
defparam \nxt_in_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt~0 (
	.dataa(!out_valid_reg1),
	.datab(!cp_ready),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt~0 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt~0 .lut_mask = 64'h1111111111111111;
defparam \nxt_uncomp_subburst_byte_cnt~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[3]~1 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!out_uncomp_byte_cnt_reg_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[3]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[3]~1 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[3]~1 .lut_mask = 64'h0FE40F4E0FE40F4E;
defparam \nxt_uncomp_subburst_byte_cnt[3]~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[4]~2 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!out_uncomp_byte_cnt_reg_2),
	.dataf(!out_uncomp_byte_cnt_reg_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[4]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[4]~2 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[4]~2 .lut_mask = 64'h00E40044FF4EFFEE;
defparam \nxt_uncomp_subburst_byte_cnt[4]~2 .shared_arith = "off";

cyclonev_lcell_comb \Add4~0 (
	.dataa(!out_uncomp_byte_cnt_reg_3),
	.datab(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datac(!out_uncomp_byte_cnt_reg_2),
	.datad(!out_uncomp_byte_cnt_reg_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add4~0 .extended_lut = "off";
defparam \Add4~0 .lut_mask = 64'h2000200020002000;
defparam \Add4~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[5]~3 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_5),
	.datae(!\Add4~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[5]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[5]~3 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[5]~3 .lut_mask = 64'h04FEAE5404FEAE54;
defparam \nxt_uncomp_subburst_byte_cnt[5]~3 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[2]~4 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[2]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[2]~4 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[2]~4 .lut_mask = 64'h0EF40EF40EF40EF4;
defparam \nxt_uncomp_subburst_byte_cnt[2]~4 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[6]~5 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_5),
	.datae(!\Add4~0_combout ),
	.dataf(!out_uncomp_byte_cnt_reg_6),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[6]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[6]~5 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[6]~5 .lut_mask = 64'h0404AE04FEFE54FE;
defparam \nxt_uncomp_subburst_byte_cnt[6]~5 .shared_arith = "off";

cyclonev_lcell_comb WideOr0(
	.dataa(!\nxt_uncomp_subburst_byte_cnt[3]~1_combout ),
	.datab(!\nxt_uncomp_subburst_byte_cnt[4]~2_combout ),
	.datac(!\nxt_uncomp_subburst_byte_cnt[5]~3_combout ),
	.datad(!\nxt_uncomp_subburst_byte_cnt[2]~4_combout ),
	.datae(!\nxt_uncomp_subburst_byte_cnt[6]~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr0.extended_lut = "off";
defparam WideOr0.lut_mask = 64'h8000000080000000;
defparam WideOr0.shared_arith = "off";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!sink0_data[69]),
	.datab(!in_ready_hold),
	.datac(!\state.ST_UNCOMP_TRANS~q ),
	.datad(!sink0_data[68]),
	.datae(!src0_valid),
	.dataf(!src0_valid1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'h0000000301010103;
defparam \Selector2~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_in_ready~3 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_in_ready~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~3 .extended_lut = "off";
defparam \nxt_in_ready~3 .lut_mask = 64'h8888888888888888;
defparam \nxt_in_ready~3 .shared_arith = "off";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!nxt_out_eop),
	.datab(!\state.ST_IDLE~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'h2222222222222222;
defparam \Selector0~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector0~1 (
	.dataa(!sink0_data[69]),
	.datab(!sink0_data[68]),
	.datac(!\state.ST_IDLE~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~1 .extended_lut = "off";
defparam \Selector0~1 .lut_mask = 64'h8080808080808080;
defparam \Selector0~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector0~2 (
	.dataa(!in_ready_hold),
	.datab(!sink0_data[68]),
	.datac(!src0_valid),
	.datad(!src_valid),
	.datae(!\Selector0~0_combout ),
	.dataf(!\Selector0~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~2 .extended_lut = "off";
defparam \Selector0~2 .lut_mask = 64'h0155FFFF0000FFFF;
defparam \Selector0~2 .shared_arith = "off";

cyclonev_lcell_comb load_next_out_cmd(
	.dataa(!out_valid_reg1),
	.datab(!cp_ready),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\load_next_out_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam load_next_out_cmd.extended_lut = "off";
defparam load_next_out_cmd.lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam load_next_out_cmd.shared_arith = "off";

dffeas \state.ST_IDLE (
	.clk(clk_clk),
	.d(\Selector0~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_IDLE~q ),
	.prn(vcc));
defparam \state.ST_IDLE .is_wysiwyg = "true";
defparam \state.ST_IDLE .power_up = "low";

cyclonev_lcell_comb \Selector2~1 (
	.dataa(!nxt_out_eop),
	.datab(!in_ready_hold),
	.datac(!\nxt_in_ready~3_combout ),
	.datad(!sink0_data[68]),
	.datae(!src0_valid),
	.dataf(!\state.ST_IDLE~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~1 .extended_lut = "off";
defparam \Selector2~1 .lut_mask = 64'h0000003300000010;
defparam \Selector2~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~2 (
	.dataa(!sink0_data[69]),
	.datab(!nxt_out_eop),
	.datac(!\nxt_in_ready~0_combout ),
	.datad(!\WideOr0~combout ),
	.datae(!\Selector2~0_combout ),
	.dataf(!\Selector2~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~2 .extended_lut = "off";
defparam \Selector2~2 .lut_mask = 64'h00C022E2AAEAAAEA;
defparam \Selector2~2 .shared_arith = "off";

dffeas \state.ST_UNCOMP_TRANS (
	.clk(clk_clk),
	.d(\Selector2~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_UNCOMP_TRANS~q ),
	.prn(vcc));
defparam \state.ST_UNCOMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_TRANS .power_up = "low";

cyclonev_lcell_comb in_valid(
	.dataa(!sink0_data[69]),
	.datab(!in_ready_hold),
	.datac(!sink0_data[68]),
	.datad(!src0_valid),
	.datae(!src0_valid1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\in_valid~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam in_valid.extended_lut = "off";
defparam in_valid.lut_mask = 64'h0003111300031113;
defparam in_valid.shared_arith = "off";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!nxt_out_eop),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'h4444444444444444;
defparam \Selector1~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~1 (
	.dataa(!sink0_data[69]),
	.datab(!stateST_COMP_TRANS),
	.datac(!nxt_out_eop),
	.datad(!\nxt_in_ready~0_combout ),
	.datae(!sink0_data[68]),
	.dataf(!\state.ST_IDLE~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~1 .extended_lut = "off";
defparam \Selector1~1 .lut_mask = 64'h8888AAAAC8CCEAEE;
defparam \Selector1~1 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[5] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[5]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[5]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[5] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[5] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[2]~4 (
	.dataa(!h2f_ARLEN_0),
	.datab(!sink0_data[69]),
	.datac(!sink0_data[68]),
	.datad(!write_cp_data_74),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[2]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[2]~4 .extended_lut = "off";
defparam \d0_int_bytes_remaining[2]~4 .lut_mask = 64'h2F222F222F222F22;
defparam \d0_int_bytes_remaining[2]~4 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[2]~5 (
	.dataa(!\new_burst_reg~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\int_bytes_remaining_reg[2]~q ),
	.datad(!\d0_int_bytes_remaining[2]~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[2]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[2]~5 .extended_lut = "off";
defparam \d0_int_bytes_remaining[2]~5 .lut_mask = 64'h287D287D287D287D;
defparam \d0_int_bytes_remaining[2]~5 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[2] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[2]~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[2]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[2] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[3]~6 (
	.dataa(!sink0_data[69]),
	.datab(!sink0_data[68]),
	.datac(!write_cp_data_75),
	.datad(!Add2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[3]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[3]~6 .extended_lut = "off";
defparam \d0_int_bytes_remaining[3]~6 .lut_mask = 64'h0357035703570357;
defparam \d0_int_bytes_remaining[3]~6 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[3]~7 (
	.dataa(!\new_burst_reg~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\int_bytes_remaining_reg[2]~q ),
	.datad(!\int_bytes_remaining_reg[3]~q ),
	.datae(!\d0_int_bytes_remaining[3]~6_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[3]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[3]~7 .extended_lut = "off";
defparam \d0_int_bytes_remaining[3]~7 .lut_mask = 64'h208A75DF208A75DF;
defparam \d0_int_bytes_remaining[3]~7 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[3] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[3]~7_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[3]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[3] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[3] .power_up = "low";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!out_byte_cnt_reg_2),
	.datab(!\int_bytes_remaining_reg[2]~q ),
	.datac(!\int_bytes_remaining_reg[3]~q ),
	.datad(!\int_bytes_remaining_reg[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'hBF40BF40BF40BF40;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[4]~8 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!sink0_data[68]),
	.datad(!\Add1~1_combout ),
	.datae(!write_cp_data_76),
	.dataf(!Add21),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[4]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[4]~8 .extended_lut = "off";
defparam \d0_int_bytes_remaining[4]~8 .lut_mask = 64'hCC00CF03DD11DF13;
defparam \d0_int_bytes_remaining[4]~8 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[4] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[4]~8_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[4]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[4] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[4] .power_up = "low";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!out_byte_cnt_reg_2),
	.datab(!\int_bytes_remaining_reg[2]~q ),
	.datac(!\int_bytes_remaining_reg[3]~q ),
	.datad(!\int_bytes_remaining_reg[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h4000400040004000;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[5]~0 (
	.dataa(!sink0_data[69]),
	.datab(!sink0_data[68]),
	.datac(!write_cp_data_77),
	.datad(!Add22),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[5]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[5]~0 .extended_lut = "off";
defparam \d0_int_bytes_remaining[5]~0 .lut_mask = 64'h0357035703570357;
defparam \d0_int_bytes_remaining[5]~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[5]~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\int_bytes_remaining_reg[5]~q ),
	.datac(!\Add1~0_combout ),
	.datad(!\d0_int_bytes_remaining[5]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[5]~1 .extended_lut = "off";
defparam \d0_int_bytes_remaining[5]~1 .lut_mask = 64'h287D287D287D287D;
defparam \d0_int_bytes_remaining[5]~1 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[6] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[6]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[6]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[6] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[6] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[6]~2 (
	.dataa(!sink0_data[69]),
	.datab(!sink0_data[68]),
	.datac(!write_cp_data_78),
	.datad(!Add23),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[6]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[6]~2 .extended_lut = "off";
defparam \d0_int_bytes_remaining[6]~2 .lut_mask = 64'h0357035703570357;
defparam \d0_int_bytes_remaining[6]~2 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[6]~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\int_bytes_remaining_reg[5]~q ),
	.datac(!\Add1~0_combout ),
	.datad(!\int_bytes_remaining_reg[6]~q ),
	.datae(!\d0_int_bytes_remaining[6]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[6]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[6]~3 .extended_lut = "off";
defparam \d0_int_bytes_remaining[6]~3 .lut_mask = 64'h08A25DF708A25DF7;
defparam \d0_int_bytes_remaining[6]~3 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!\d0_int_bytes_remaining[2]~5_combout ),
	.datab(!\d0_int_bytes_remaining[3]~7_combout ),
	.datac(!\d0_int_bytes_remaining[4]~8_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'h4040404040404040;
defparam \Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \new_burst_reg~0 (
	.dataa(!\in_valid~combout ),
	.datab(!\Selector1~0_combout ),
	.datac(!\Selector1~1_combout ),
	.datad(!\d0_int_bytes_remaining[5]~1_combout ),
	.datae(!\d0_int_bytes_remaining[6]~3_combout ),
	.dataf(!\Equal0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\new_burst_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \new_burst_reg~0 .extended_lut = "off";
defparam \new_burst_reg~0 .lut_mask = 64'h8C8C8C8CFF8C8C8C;
defparam \new_burst_reg~0 .shared_arith = "off";

dffeas new_burst_reg(
	.clk(clk_clk),
	.d(\new_burst_reg~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\new_burst_reg~q ),
	.prn(vcc));
defparam new_burst_reg.is_wysiwyg = "true";
defparam new_burst_reg.power_up = "low";

cyclonev_lcell_comb \Selector1~2 (
	.dataa(!in_ready_hold),
	.datab(!sink0_data[68]),
	.datac(!src0_valid),
	.datad(!src_valid),
	.datae(!\Selector1~0_combout ),
	.dataf(!\Selector1~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~2 .extended_lut = "off";
defparam \Selector1~2 .lut_mask = 64'h0155FFFF0000FFFF;
defparam \Selector1~2 .shared_arith = "off";

cyclonev_lcell_comb \WideNor0~1 (
	.dataa(!sink0_data[69]),
	.datab(!sink0_data[68]),
	.datac(!WideNor0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideNor0~1 .extended_lut = "off";
defparam \WideNor0~1 .lut_mask = 64'h8A8A8A8A8A8A8A8A;
defparam \WideNor0~1 .shared_arith = "off";

cyclonev_lcell_comb \NON_PIPELINED_INPUTS.load_next_cmd (
	.dataa(!in_ready_hold),
	.datab(!nxt_in_ready1),
	.datac(!nxt_in_ready),
	.datad(!sink0_data[68]),
	.datae(!src0_valid),
	.dataf(!src_valid),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \NON_PIPELINED_INPUTS.load_next_cmd .extended_lut = "off";
defparam \NON_PIPELINED_INPUTS.load_next_cmd .lut_mask = 64'h0000001515151515;
defparam \NON_PIPELINED_INPUTS.load_next_cmd .shared_arith = "off";

dffeas in_bytecount_reg_zero(
	.clk(clk_clk),
	.d(\WideNor0~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_bytecount_reg_zero~q ),
	.prn(vcc));
defparam in_bytecount_reg_zero.is_wysiwyg = "true";
defparam in_bytecount_reg_zero.power_up = "low";

cyclonev_lcell_comb \nxt_out_valid~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!\new_burst_reg~q ),
	.datac(!mem_used_1),
	.datad(!\in_bytecount_reg_zero~q ),
	.datae(!cp_ready1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_valid~0 .extended_lut = "off";
defparam \nxt_out_valid~0 .lut_mask = 64'h4540550045405500;
defparam \nxt_out_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_out_valid~1 (
	.dataa(!in_ready_hold),
	.datab(!sink0_data[68]),
	.datac(!src0_valid),
	.datad(!src_valid),
	.datae(!\nxt_out_valid~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_valid~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_valid~1 .extended_lut = "off";
defparam \nxt_out_valid~1 .lut_mask = 64'h0155FFFF0155FFFF;
defparam \nxt_out_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!sink0_data[87]),
	.datab(!sink0_data[88]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h8888888888888888;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~0 (
	.dataa(!nxt_out_eop),
	.datab(!\nxt_in_ready~0_combout ),
	.datac(!\WideOr0~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'h8080808080808080;
defparam \Selector3~0 .shared_arith = "off";

dffeas \in_size_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[86]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[0]~q ),
	.prn(vcc));
defparam \in_size_reg[0] .is_wysiwyg = "true";
defparam \in_size_reg[0] .power_up = "low";

dffeas \in_size_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[87]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[1]~q ),
	.prn(vcc));
defparam \in_size_reg[1] .is_wysiwyg = "true";
defparam \in_size_reg[1] .power_up = "low";

dffeas \in_size_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[88]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[2]~q ),
	.prn(vcc));
defparam \in_size_reg[2] .is_wysiwyg = "true";
defparam \in_size_reg[2] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[87]),
	.datac(!sink0_data[88]),
	.datad(!\in_size_reg[1]~q ),
	.datae(!\in_size_reg[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~0 .extended_lut = "off";
defparam \ShiftLeft0~0 .lut_mask = 64'h10BA101010BA1010;
defparam \ShiftLeft0~0 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~1 .extended_lut = "off";
defparam \ShiftLeft0~1 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~1 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[3] (
	.clk(clk_clk),
	.d(\ShiftLeft0~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[3]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[3] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[3] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~2 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~2 .extended_lut = "off";
defparam \ShiftLeft0~2 .lut_mask = 64'h00E400E400E400E4;
defparam \ShiftLeft0~2 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[2] (
	.clk(clk_clk),
	.d(\ShiftLeft0~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[2]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[2] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[2] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[87]),
	.datac(!sink0_data[88]),
	.datad(!\in_size_reg[1]~q ),
	.datae(!\in_size_reg[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~3 .extended_lut = "off";
defparam \ShiftLeft0~3 .lut_mask = 64'hEA404040EA404040;
defparam \ShiftLeft0~3 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~4 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~4 .extended_lut = "off";
defparam \ShiftLeft0~4 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~4 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[1] (
	.clk(clk_clk),
	.d(\ShiftLeft0~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[1]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[1] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[1] .power_up = "low";

dffeas \int_byte_cnt_narrow_reg[0] (
	.clk(clk_clk),
	.d(\align_address_to_size|LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[0]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[0] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[0] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[0]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~3 (
	.dataa(!h2f_ARADDR_0),
	.datab(!sink0_data[69]),
	.datac(!sink0_data[68]),
	.datad(!out_data_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~3 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~3 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[0]~3 .shared_arith = "off";

dffeas \in_burstwrap_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[79]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[0]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[0] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[0] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[0]~0 (
	.dataa(!Selector13),
	.datab(!Selector6),
	.datac(!sink0_data[68]),
	.datad(!sink0_data[69]),
	.datae(!\new_burst_reg~q ),
	.dataf(!\d0_int_nxt_addr[0]~4_combout ),
	.datag(!\in_burstwrap_reg[0]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[0]~0 .extended_lut = "on";
defparam \nxt_addr[0]~0 .lut_mask = 64'h00000000F0F0FCA8;
defparam \nxt_addr[0]~0 .shared_arith = "off";

dffeas \int_nxt_addr_reg[0] (
	.clk(clk_clk),
	.d(\nxt_addr[0]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[0] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~4 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\Add0~13_sumout ),
	.datac(!\align_address_to_size|LessThan0~0_combout ),
	.datad(!\d0_int_nxt_addr[0]~3_combout ),
	.datae(!\int_nxt_addr_reg[0]~q ),
	.dataf(!\in_burstwrap_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~4 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~4 .lut_mask = 64'h0005AAAF2227AAAF;
defparam \d0_int_nxt_addr[0]~4 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[0] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[0]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[0] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[1]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[1]~q ),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \in_burstwrap_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[80]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[1]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[1] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[1] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[1]~4 (
	.dataa(!Selector12),
	.datab(!Selector5),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!\new_burst_reg~q ),
	.dataf(!\d0_int_nxt_addr[1]~2_combout ),
	.datag(!\in_burstwrap_reg[1]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[1]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[1]~4 .extended_lut = "on";
defparam \nxt_addr[1]~4 .lut_mask = 64'h00000000F0F0FAC8;
defparam \nxt_addr[1]~4 .shared_arith = "off";

dffeas \int_nxt_addr_reg[1] (
	.clk(clk_clk),
	.d(\nxt_addr[1]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[1] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~7 (
	.dataa(!h2f_ARADDR_1),
	.datab(!sink0_data[69]),
	.datac(!sink0_data[68]),
	.datad(!out_data_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~7 .extended_lut = "off";
defparam \d0_int_nxt_addr[1]~7 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[1]~7 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~2 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\Add0~9_sumout ),
	.datac(!\in_burstwrap_reg[1]~q ),
	.datad(!\int_nxt_addr_reg[1]~q ),
	.datae(!\ShiftLeft0~3_combout ),
	.dataf(!\d0_int_nxt_addr[1]~7_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~2 .extended_lut = "off";
defparam \d0_int_nxt_addr[1]~2 .lut_mask = 64'h02AA02AA02AA57FF;
defparam \d0_int_nxt_addr[1]~2 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[1] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[1]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[1] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_2),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[2]~q ),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[3]~q ),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

dffeas \in_burstwrap_reg[3] (
	.clk(clk_clk),
	.d(sink0_data[82]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[3]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[3] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[3] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[3]~12 (
	.dataa(!Selector10),
	.datab(!Selector3),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!\new_burst_reg~q ),
	.dataf(!\d0_int_nxt_addr[3]~0_combout ),
	.datag(!\in_burstwrap_reg[3]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[3]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[3]~12 .extended_lut = "on";
defparam \nxt_addr[3]~12 .lut_mask = 64'h00000000F0F0FAC8;
defparam \nxt_addr[3]~12 .shared_arith = "off";

dffeas \int_nxt_addr_reg[3] (
	.clk(clk_clk),
	.d(\nxt_addr[3]~12_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[3]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[3] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~5 (
	.dataa(!\Add0~1_sumout ),
	.datab(!\in_burstwrap_reg[3]~q ),
	.datac(!\int_nxt_addr_reg[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~5 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~5 .lut_mask = 64'hE0E0E0E0E0E0E0E0;
defparam \d0_int_nxt_addr[3]~5 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!h2f_ARADDR_3),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!base_address_3),
	.dataf(!\d0_int_nxt_addr[3]~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~0 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~0 .lut_mask = 64'hABABABFF01010155;
defparam \d0_int_nxt_addr[3]~0 .shared_arith = "off";

dffeas \in_burstwrap_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[81]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[2]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[2] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[2] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[2]~8 (
	.dataa(!Selector11),
	.datab(!Selector4),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!\new_burst_reg~q ),
	.dataf(!\d0_int_nxt_addr[2]~1_combout ),
	.datag(!\in_burstwrap_reg[2]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[2]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[2]~8 .extended_lut = "on";
defparam \nxt_addr[2]~8 .lut_mask = 64'h00000000F0F0FAC8;
defparam \nxt_addr[2]~8 .shared_arith = "off";

dffeas \int_nxt_addr_reg[2] (
	.clk(clk_clk),
	.d(\nxt_addr[2]~8_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[2]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~6 (
	.dataa(!\Add0~5_sumout ),
	.datab(!\in_burstwrap_reg[2]~q ),
	.datac(!\int_nxt_addr_reg[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~6 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~6 .lut_mask = 64'hE0E0E0E0E0E0E0E0;
defparam \d0_int_nxt_addr[2]~6 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!h2f_ARADDR_2),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!base_address_2),
	.dataf(!\d0_int_nxt_addr[2]~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~1 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~1 .lut_mask = 64'hABABABFF01010155;
defparam \d0_int_nxt_addr[2]~1 .shared_arith = "off";

dffeas in_eop_reg(
	.clk(clk_clk),
	.d(sink0_endofpacket),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_eop_reg~q ),
	.prn(vcc));
defparam in_eop_reg.is_wysiwyg = "true";
defparam in_eop_reg.power_up = "low";

endmodule

module spw_babasu_altera_merlin_address_alignment_7 (
	new_burst_reg,
	src_data_86,
	in_size_reg_0,
	ShiftLeft0,
	LessThan0)/* synthesis synthesis_greybox=0 */;
input 	new_burst_reg;
input 	src_data_86;
input 	in_size_reg_0;
input 	ShiftLeft0;
output 	LessThan0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!new_burst_reg),
	.datab(!src_data_86),
	.datac(!in_size_reg_0),
	.datad(!ShiftLeft0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan0),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h00E400E400E400E4;
defparam \LessThan0~0 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_burst_adapter_7 (
	h2f_ARADDR_0,
	h2f_ARADDR_1,
	h2f_ARADDR_2,
	h2f_ARADDR_3,
	h2f_ARLEN_0,
	nxt_in_ready,
	in_ready_hold,
	stateST_COMP_TRANS,
	out_valid_reg,
	in_narrow_reg,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	in_data_reg_68,
	cp_ready,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready1,
	saved_grant_1,
	Equal9,
	saved_grant_0,
	altera_reset_synchronizer_int_chain_out,
	in_data_reg_0,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	Add2,
	Add21,
	Add22,
	Add23,
	Equal5,
	write_cp_data_77,
	write_cp_data_78,
	write_cp_data_75,
	write_cp_data_74,
	write_cp_data_76,
	WideNor0,
	nxt_out_eop,
	src9_valid,
	src_valid,
	cp_ready1,
	in_data_reg_69,
	src_data_87,
	src_data_88,
	src_valid1,
	src_data_35,
	src_data_34,
	src_data_33,
	src_data_32,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_6,
	src_payload_0,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	Selector3,
	Selector10,
	base_address_3,
	Selector4,
	Selector11,
	base_address_2,
	src_payload,
	src_data_82,
	src_data_81,
	src_data_105,
	src_data_106,
	src_data_107,
	src_data_108,
	src_data_109,
	src_data_110,
	src_data_111,
	src_data_112,
	src_data_113,
	src_data_114,
	src_data_115,
	src_data_116,
	src_data_86,
	Selector5,
	Selector12,
	out_data_1,
	src_data_80,
	out_data_0,
	Selector6,
	Selector13,
	src_data_79,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARADDR_0;
input 	h2f_ARADDR_1;
input 	h2f_ARADDR_2;
input 	h2f_ARADDR_3;
input 	h2f_ARLEN_0;
output 	nxt_in_ready;
input 	in_ready_hold;
output 	stateST_COMP_TRANS;
output 	out_valid_reg;
output 	in_narrow_reg;
output 	in_byteen_reg_3;
output 	in_byteen_reg_2;
output 	in_byteen_reg_1;
output 	in_byteen_reg_0;
output 	in_data_reg_68;
input 	cp_ready;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready1;
input 	saved_grant_1;
input 	Equal9;
input 	saved_grant_0;
input 	altera_reset_synchronizer_int_chain_out;
output 	in_data_reg_0;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
input 	Add2;
input 	Add21;
input 	Add22;
input 	Add23;
input 	Equal5;
input 	write_cp_data_77;
input 	write_cp_data_78;
input 	write_cp_data_75;
input 	write_cp_data_74;
input 	write_cp_data_76;
input 	WideNor0;
output 	nxt_out_eop;
input 	src9_valid;
input 	src_valid;
input 	cp_ready1;
output 	in_data_reg_69;
input 	src_data_87;
input 	src_data_88;
input 	src_valid1;
input 	src_data_35;
input 	src_data_34;
input 	src_data_33;
input 	src_data_32;
output 	out_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_6;
input 	src_payload_0;
output 	in_data_reg_105;
output 	in_data_reg_106;
output 	in_data_reg_107;
output 	in_data_reg_108;
output 	in_data_reg_109;
output 	in_data_reg_110;
output 	in_data_reg_111;
output 	in_data_reg_112;
output 	in_data_reg_113;
output 	in_data_reg_114;
output 	in_data_reg_115;
output 	in_data_reg_116;
input 	Selector3;
input 	Selector10;
input 	base_address_3;
input 	Selector4;
input 	Selector11;
input 	base_address_2;
input 	src_payload;
input 	src_data_82;
input 	src_data_81;
input 	src_data_105;
input 	src_data_106;
input 	src_data_107;
input 	src_data_108;
input 	src_data_109;
input 	src_data_110;
input 	src_data_111;
input 	src_data_112;
input 	src_data_113;
input 	src_data_114;
input 	src_data_115;
input 	src_data_116;
input 	src_data_86;
input 	Selector5;
input 	Selector12;
input 	out_data_1;
input 	src_data_80;
input 	out_data_0;
input 	Selector6;
input 	Selector13;
input 	src_data_79;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



spw_babasu_altera_merlin_burst_adapter_13_1_7 \altera_merlin_burst_adapter_13_1.burst_adapter (
	.h2f_ARADDR_0(h2f_ARADDR_0),
	.h2f_ARADDR_1(h2f_ARADDR_1),
	.h2f_ARADDR_2(h2f_ARADDR_2),
	.h2f_ARADDR_3(h2f_ARADDR_3),
	.h2f_ARLEN_0(h2f_ARLEN_0),
	.nxt_in_ready(nxt_in_ready),
	.in_ready_hold(in_ready_hold),
	.stateST_COMP_TRANS(stateST_COMP_TRANS),
	.out_valid_reg1(out_valid_reg),
	.in_narrow_reg1(in_narrow_reg),
	.in_byteen_reg_3(in_byteen_reg_3),
	.in_byteen_reg_2(in_byteen_reg_2),
	.in_byteen_reg_1(in_byteen_reg_1),
	.in_byteen_reg_0(in_byteen_reg_0),
	.in_data_reg_68(in_data_reg_68),
	.cp_ready(cp_ready),
	.stateST_UNCOMP_WR_SUBBURST(stateST_UNCOMP_WR_SUBBURST),
	.nxt_in_ready1(nxt_in_ready1),
	.sink0_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_116,src_data_115,src_data_114,src_data_113,src_data_112,src_data_111,src_data_110,src_data_109,src_data_108,src_data_107,src_data_106,src_data_105,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_88,src_data_87,
src_data_86,gnd,gnd,gnd,src_data_82,src_data_81,src_data_80,src_data_79,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,saved_grant_1,saved_grant_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_35,src_data_34,src_data_33,
src_data_32,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_payload}),
	.Equal9(Equal9),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.in_data_reg_0(in_data_reg_0),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_3),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_2),
	.Add2(Add2),
	.Add21(Add21),
	.Add22(Add22),
	.Add23(Add23),
	.Equal5(Equal5),
	.write_cp_data_77(write_cp_data_77),
	.write_cp_data_78(write_cp_data_78),
	.write_cp_data_75(write_cp_data_75),
	.write_cp_data_74(write_cp_data_74),
	.write_cp_data_76(write_cp_data_76),
	.WideNor0(WideNor0),
	.nxt_out_eop(nxt_out_eop),
	.src9_valid(src9_valid),
	.src_valid(src_valid),
	.cp_ready1(cp_ready1),
	.in_data_reg_69(in_data_reg_69),
	.src_valid1(src_valid1),
	.out_byte_cnt_reg_2(out_byte_cnt_reg_2),
	.out_uncomp_byte_cnt_reg_4(out_uncomp_byte_cnt_reg_4),
	.out_uncomp_byte_cnt_reg_3(out_uncomp_byte_cnt_reg_3),
	.out_uncomp_byte_cnt_reg_2(out_uncomp_byte_cnt_reg_2),
	.out_uncomp_byte_cnt_reg_5(out_uncomp_byte_cnt_reg_5),
	.out_uncomp_byte_cnt_reg_6(out_uncomp_byte_cnt_reg_6),
	.sink0_endofpacket(src_payload_0),
	.in_data_reg_105(in_data_reg_105),
	.in_data_reg_106(in_data_reg_106),
	.in_data_reg_107(in_data_reg_107),
	.in_data_reg_108(in_data_reg_108),
	.in_data_reg_109(in_data_reg_109),
	.in_data_reg_110(in_data_reg_110),
	.in_data_reg_111(in_data_reg_111),
	.in_data_reg_112(in_data_reg_112),
	.in_data_reg_113(in_data_reg_113),
	.in_data_reg_114(in_data_reg_114),
	.in_data_reg_115(in_data_reg_115),
	.in_data_reg_116(in_data_reg_116),
	.Selector3(Selector3),
	.Selector10(Selector10),
	.base_address_3(base_address_3),
	.Selector4(Selector4),
	.Selector11(Selector11),
	.base_address_2(base_address_2),
	.Selector5(Selector5),
	.Selector12(Selector12),
	.out_data_1(out_data_1),
	.out_data_0(out_data_0),
	.Selector6(Selector6),
	.Selector13(Selector13),
	.clk_clk(clk_clk));

endmodule

module spw_babasu_altera_merlin_burst_adapter_13_1_7 (
	h2f_ARADDR_0,
	h2f_ARADDR_1,
	h2f_ARADDR_2,
	h2f_ARADDR_3,
	h2f_ARLEN_0,
	nxt_in_ready,
	in_ready_hold,
	stateST_COMP_TRANS,
	out_valid_reg1,
	in_narrow_reg1,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	in_data_reg_68,
	cp_ready,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready1,
	sink0_data,
	Equal9,
	altera_reset_synchronizer_int_chain_out,
	in_data_reg_0,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	Add2,
	Add21,
	Add22,
	Add23,
	Equal5,
	write_cp_data_77,
	write_cp_data_78,
	write_cp_data_75,
	write_cp_data_74,
	write_cp_data_76,
	WideNor0,
	nxt_out_eop,
	src9_valid,
	src_valid,
	cp_ready1,
	in_data_reg_69,
	src_valid1,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_6,
	sink0_endofpacket,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	Selector3,
	Selector10,
	base_address_3,
	Selector4,
	Selector11,
	base_address_2,
	Selector5,
	Selector12,
	out_data_1,
	out_data_0,
	Selector6,
	Selector13,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARADDR_0;
input 	h2f_ARADDR_1;
input 	h2f_ARADDR_2;
input 	h2f_ARADDR_3;
input 	h2f_ARLEN_0;
output 	nxt_in_ready;
input 	in_ready_hold;
output 	stateST_COMP_TRANS;
output 	out_valid_reg1;
output 	in_narrow_reg1;
output 	in_byteen_reg_3;
output 	in_byteen_reg_2;
output 	in_byteen_reg_1;
output 	in_byteen_reg_0;
output 	in_data_reg_68;
input 	cp_ready;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready1;
input 	[128:0] sink0_data;
input 	Equal9;
input 	altera_reset_synchronizer_int_chain_out;
output 	in_data_reg_0;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
input 	Add2;
input 	Add21;
input 	Add22;
input 	Add23;
input 	Equal5;
input 	write_cp_data_77;
input 	write_cp_data_78;
input 	write_cp_data_75;
input 	write_cp_data_74;
input 	write_cp_data_76;
input 	WideNor0;
output 	nxt_out_eop;
input 	src9_valid;
input 	src_valid;
input 	cp_ready1;
output 	in_data_reg_69;
input 	src_valid1;
output 	out_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_6;
input 	sink0_endofpacket;
output 	in_data_reg_105;
output 	in_data_reg_106;
output 	in_data_reg_107;
output 	in_data_reg_108;
output 	in_data_reg_109;
output 	in_data_reg_110;
output 	in_data_reg_111;
output 	in_data_reg_112;
output 	in_data_reg_113;
output 	in_data_reg_114;
output 	in_data_reg_115;
output 	in_data_reg_116;
input 	Selector3;
input 	Selector10;
input 	base_address_3;
input 	Selector4;
input 	Selector11;
input 	base_address_2;
input 	Selector5;
input 	Selector12;
input 	out_data_1;
input 	out_data_0;
input 	Selector6;
input 	Selector13;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \align_address_to_size|LessThan0~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt[4]~1_combout ;
wire \nxt_uncomp_subburst_byte_cnt[3]~2_combout ;
wire \Add4~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt[5]~3_combout ;
wire \nxt_uncomp_subburst_byte_cnt[2]~4_combout ;
wire \nxt_uncomp_subburst_byte_cnt[6]~5_combout ;
wire \WideOr0~combout ;
wire \in_valid~combout ;
wire \Selector0~0_combout ;
wire \load_next_out_cmd~combout ;
wire \state.ST_IDLE~q ;
wire \Selector2~0_combout ;
wire \Selector2~1_combout ;
wire \Selector2~2_combout ;
wire \state.ST_UNCOMP_TRANS~q ;
wire \Selector1~0_combout ;
wire \Selector1~1_combout ;
wire \int_bytes_remaining_reg[3]~q ;
wire \d0_int_bytes_remaining[2]~2_combout ;
wire \d0_int_bytes_remaining[2]~3_combout ;
wire \int_bytes_remaining_reg[2]~q ;
wire \d0_int_bytes_remaining[3]~0_combout ;
wire \d0_int_bytes_remaining[3]~1_combout ;
wire \int_bytes_remaining_reg[6]~q ;
wire \Add1~1_combout ;
wire \d0_int_bytes_remaining[4]~8_combout ;
wire \int_bytes_remaining_reg[4]~q ;
wire \Add1~0_combout ;
wire \d0_int_bytes_remaining[5]~6_combout ;
wire \d0_int_bytes_remaining[5]~7_combout ;
wire \int_bytes_remaining_reg[5]~q ;
wire \d0_int_bytes_remaining[6]~4_combout ;
wire \d0_int_bytes_remaining[6]~5_combout ;
wire \new_burst_reg~0_combout ;
wire \new_burst_reg~q ;
wire \WideNor0~0_combout ;
wire \NON_PIPELINED_INPUTS.load_next_cmd~combout ;
wire \in_bytecount_reg_zero~q ;
wire \nxt_out_valid~0_combout ;
wire \LessThan0~0_combout ;
wire \Selector3~0_combout ;
wire \in_size_reg[0]~q ;
wire \in_size_reg[1]~q ;
wire \in_size_reg[2]~q ;
wire \ShiftLeft0~0_combout ;
wire \ShiftLeft0~1_combout ;
wire \int_byte_cnt_narrow_reg[3]~q ;
wire \ShiftLeft0~2_combout ;
wire \int_byte_cnt_narrow_reg[2]~q ;
wire \ShiftLeft0~3_combout ;
wire \ShiftLeft0~4_combout ;
wire \int_byte_cnt_narrow_reg[1]~q ;
wire \int_byte_cnt_narrow_reg[0]~q ;
wire \Add0~13_sumout ;
wire \d0_int_nxt_addr[0]~3_combout ;
wire \in_burstwrap_reg[0]~q ;
wire \nxt_addr[0]~0_combout ;
wire \int_nxt_addr_reg[0]~q ;
wire \d0_int_nxt_addr[0]~4_combout ;
wire \int_nxt_addr_reg_dly[0]~q ;
wire \Add0~14 ;
wire \Add0~9_sumout ;
wire \in_burstwrap_reg[1]~q ;
wire \nxt_addr[1]~4_combout ;
wire \int_nxt_addr_reg[1]~q ;
wire \d0_int_nxt_addr[1]~7_combout ;
wire \d0_int_nxt_addr[1]~2_combout ;
wire \int_nxt_addr_reg_dly[1]~q ;
wire \Add0~10 ;
wire \Add0~6 ;
wire \Add0~1_sumout ;
wire \in_burstwrap_reg[3]~q ;
wire \nxt_addr[3]~12_combout ;
wire \int_nxt_addr_reg[3]~q ;
wire \d0_int_nxt_addr[3]~5_combout ;
wire \d0_int_nxt_addr[3]~0_combout ;
wire \Add0~5_sumout ;
wire \in_burstwrap_reg[2]~q ;
wire \nxt_addr[2]~8_combout ;
wire \int_nxt_addr_reg[2]~q ;
wire \d0_int_nxt_addr[2]~6_combout ;
wire \d0_int_nxt_addr[2]~1_combout ;
wire \in_eop_reg~q ;


spw_babasu_altera_merlin_address_alignment_8 align_address_to_size(
	.new_burst_reg(\new_burst_reg~q ),
	.src_data_86(sink0_data[86]),
	.in_size_reg_0(\in_size_reg[0]~q ),
	.ShiftLeft0(\ShiftLeft0~3_combout ),
	.LessThan0(\align_address_to_size|LessThan0~0_combout ));

cyclonev_lcell_comb \nxt_in_ready~1 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!in_ready_hold),
	.datac(!out_valid_reg1),
	.datad(!cp_ready),
	.datae(!stateST_COMP_TRANS),
	.dataf(!\new_burst_reg~q ),
	.datag(!stateST_UNCOMP_WR_SUBBURST),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~1 .extended_lut = "on";
defparam \nxt_in_ready~1 .lut_mask = 64'h2020F0F02020F0FF;
defparam \nxt_in_ready~1 .shared_arith = "off";

dffeas \state.ST_COMP_TRANS (
	.clk(clk_clk),
	.d(\Selector1~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_COMP_TRANS),
	.prn(vcc));
defparam \state.ST_COMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_COMP_TRANS .power_up = "low";

dffeas out_valid_reg(
	.clk(clk_clk),
	.d(\nxt_out_valid~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_valid_reg1),
	.prn(vcc));
defparam out_valid_reg.is_wysiwyg = "true";
defparam out_valid_reg.power_up = "low";

dffeas in_narrow_reg(
	.clk(clk_clk),
	.d(\LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_narrow_reg1),
	.prn(vcc));
defparam in_narrow_reg.is_wysiwyg = "true";
defparam in_narrow_reg.power_up = "low";

dffeas \in_byteen_reg[3] (
	.clk(clk_clk),
	.d(sink0_data[35]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_3),
	.prn(vcc));
defparam \in_byteen_reg[3] .is_wysiwyg = "true";
defparam \in_byteen_reg[3] .power_up = "low";

dffeas \in_byteen_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[34]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_2),
	.prn(vcc));
defparam \in_byteen_reg[2] .is_wysiwyg = "true";
defparam \in_byteen_reg[2] .power_up = "low";

dffeas \in_byteen_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[33]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_1),
	.prn(vcc));
defparam \in_byteen_reg[1] .is_wysiwyg = "true";
defparam \in_byteen_reg[1] .power_up = "low";

dffeas \in_byteen_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[32]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_0),
	.prn(vcc));
defparam \in_byteen_reg[0] .is_wysiwyg = "true";
defparam \in_byteen_reg[0] .power_up = "low";

dffeas \in_data_reg[68] (
	.clk(clk_clk),
	.d(sink0_data[68]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_68),
	.prn(vcc));
defparam \in_data_reg[68] .is_wysiwyg = "true";
defparam \in_data_reg[68] .power_up = "low";

dffeas \state.ST_UNCOMP_WR_SUBBURST (
	.clk(clk_clk),
	.d(\Selector3~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_UNCOMP_WR_SUBBURST),
	.prn(vcc));
defparam \state.ST_UNCOMP_WR_SUBBURST .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_WR_SUBBURST .power_up = "low";

cyclonev_lcell_comb \nxt_in_ready~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!out_valid_reg1),
	.datac(!cp_ready),
	.datad(!\state.ST_UNCOMP_TRANS~q ),
	.datae(!stateST_UNCOMP_WR_SUBBURST),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~0 .extended_lut = "off";
defparam \nxt_in_ready~0 .lut_mask = 64'h008A8A8A008A8A8A;
defparam \nxt_in_ready~0 .shared_arith = "off";

dffeas \in_data_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[0]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_0),
	.prn(vcc));
defparam \in_data_reg[0] .is_wysiwyg = "true";
defparam \in_data_reg[0] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[3] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[3]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_3),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[3] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[2] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[2]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_2),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[2] .power_up = "low";

cyclonev_lcell_comb \nxt_out_eop~0 (
	.dataa(!\in_eop_reg~q ),
	.datab(!stateST_COMP_TRANS),
	.datac(!\new_burst_reg~q ),
	.datad(!cp_ready),
	.datae(!\in_bytecount_reg_zero~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_out_eop),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_eop~0 .extended_lut = "off";
defparam \nxt_out_eop~0 .lut_mask = 64'h4447774744477747;
defparam \nxt_out_eop~0 .shared_arith = "off";

dffeas \in_data_reg[69] (
	.clk(clk_clk),
	.d(sink0_data[69]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_69),
	.prn(vcc));
defparam \in_data_reg[69] .is_wysiwyg = "true";
defparam \in_data_reg[69] .power_up = "low";

dffeas \out_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[4] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[4]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_4),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[4] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[4] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[3] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[3]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_3),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[3] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[3] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[2]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[5] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[5]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_5),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[5] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[5] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[6] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[6]~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_6),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[6] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[6] .power_up = "low";

dffeas \in_data_reg[105] (
	.clk(clk_clk),
	.d(sink0_data[105]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_105),
	.prn(vcc));
defparam \in_data_reg[105] .is_wysiwyg = "true";
defparam \in_data_reg[105] .power_up = "low";

dffeas \in_data_reg[106] (
	.clk(clk_clk),
	.d(sink0_data[106]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_106),
	.prn(vcc));
defparam \in_data_reg[106] .is_wysiwyg = "true";
defparam \in_data_reg[106] .power_up = "low";

dffeas \in_data_reg[107] (
	.clk(clk_clk),
	.d(sink0_data[107]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_107),
	.prn(vcc));
defparam \in_data_reg[107] .is_wysiwyg = "true";
defparam \in_data_reg[107] .power_up = "low";

dffeas \in_data_reg[108] (
	.clk(clk_clk),
	.d(sink0_data[108]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_108),
	.prn(vcc));
defparam \in_data_reg[108] .is_wysiwyg = "true";
defparam \in_data_reg[108] .power_up = "low";

dffeas \in_data_reg[109] (
	.clk(clk_clk),
	.d(sink0_data[109]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_109),
	.prn(vcc));
defparam \in_data_reg[109] .is_wysiwyg = "true";
defparam \in_data_reg[109] .power_up = "low";

dffeas \in_data_reg[110] (
	.clk(clk_clk),
	.d(sink0_data[110]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_110),
	.prn(vcc));
defparam \in_data_reg[110] .is_wysiwyg = "true";
defparam \in_data_reg[110] .power_up = "low";

dffeas \in_data_reg[111] (
	.clk(clk_clk),
	.d(sink0_data[111]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_111),
	.prn(vcc));
defparam \in_data_reg[111] .is_wysiwyg = "true";
defparam \in_data_reg[111] .power_up = "low";

dffeas \in_data_reg[112] (
	.clk(clk_clk),
	.d(sink0_data[112]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_112),
	.prn(vcc));
defparam \in_data_reg[112] .is_wysiwyg = "true";
defparam \in_data_reg[112] .power_up = "low";

dffeas \in_data_reg[113] (
	.clk(clk_clk),
	.d(sink0_data[113]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_113),
	.prn(vcc));
defparam \in_data_reg[113] .is_wysiwyg = "true";
defparam \in_data_reg[113] .power_up = "low";

dffeas \in_data_reg[114] (
	.clk(clk_clk),
	.d(sink0_data[114]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_114),
	.prn(vcc));
defparam \in_data_reg[114] .is_wysiwyg = "true";
defparam \in_data_reg[114] .power_up = "low";

dffeas \in_data_reg[115] (
	.clk(clk_clk),
	.d(sink0_data[115]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_115),
	.prn(vcc));
defparam \in_data_reg[115] .is_wysiwyg = "true";
defparam \in_data_reg[115] .power_up = "low";

dffeas \in_data_reg[116] (
	.clk(clk_clk),
	.d(sink0_data[116]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_116),
	.prn(vcc));
defparam \in_data_reg[116] .is_wysiwyg = "true";
defparam \in_data_reg[116] .power_up = "low";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt~0 (
	.dataa(!out_valid_reg1),
	.datab(!cp_ready),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt~0 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt~0 .lut_mask = 64'h1111111111111111;
defparam \nxt_uncomp_subburst_byte_cnt~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[4]~1 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!out_uncomp_byte_cnt_reg_3),
	.datae(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.dataf(!out_uncomp_byte_cnt_reg_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[4]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[4]~1 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[4]~1 .lut_mask = 64'h0F0FE44E0F0F4E4E;
defparam \nxt_uncomp_subburst_byte_cnt[4]~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[3]~2 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!out_uncomp_byte_cnt_reg_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[3]~2 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[3]~2 .lut_mask = 64'h0FE40F4E0FE40F4E;
defparam \nxt_uncomp_subburst_byte_cnt[3]~2 .shared_arith = "off";

cyclonev_lcell_comb \Add4~0 (
	.dataa(!out_uncomp_byte_cnt_reg_4),
	.datab(!out_uncomp_byte_cnt_reg_3),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add4~0 .extended_lut = "off";
defparam \Add4~0 .lut_mask = 64'h0800080008000800;
defparam \Add4~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[5]~3 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_5),
	.datae(!\Add4~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[5]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[5]~3 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[5]~3 .lut_mask = 64'h04FEAE5404FEAE54;
defparam \nxt_uncomp_subburst_byte_cnt[5]~3 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[2]~4 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[2]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[2]~4 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[2]~4 .lut_mask = 64'h0EF40EF40EF40EF4;
defparam \nxt_uncomp_subburst_byte_cnt[2]~4 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[6]~5 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_5),
	.datae(!\Add4~0_combout ),
	.dataf(!out_uncomp_byte_cnt_reg_6),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[6]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[6]~5 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[6]~5 .lut_mask = 64'h0404AE04FEFE54FE;
defparam \nxt_uncomp_subburst_byte_cnt[6]~5 .shared_arith = "off";

cyclonev_lcell_comb WideOr0(
	.dataa(!\nxt_uncomp_subburst_byte_cnt[4]~1_combout ),
	.datab(!\nxt_uncomp_subburst_byte_cnt[3]~2_combout ),
	.datac(!\nxt_uncomp_subburst_byte_cnt[5]~3_combout ),
	.datad(!\nxt_uncomp_subburst_byte_cnt[2]~4_combout ),
	.datae(!\nxt_uncomp_subburst_byte_cnt[6]~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr0.extended_lut = "off";
defparam WideOr0.lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam WideOr0.shared_arith = "off";

cyclonev_lcell_comb in_valid(
	.dataa(!in_ready_hold),
	.datab(!Equal5),
	.datac(!Equal9),
	.datad(!sink0_data[68]),
	.datae(!src9_valid),
	.dataf(!src_valid),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\in_valid~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam in_valid.extended_lut = "off";
defparam in_valid.lut_mask = 64'h0000000155555555;
defparam in_valid.shared_arith = "off";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!sink0_data[69]),
	.datab(!nxt_out_eop),
	.datac(!sink0_data[68]),
	.datad(!\in_valid~combout ),
	.datae(!\state.ST_IDLE~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'h005FCCFF005FCCFF;
defparam \Selector0~0 .shared_arith = "off";

cyclonev_lcell_comb load_next_out_cmd(
	.dataa(!out_valid_reg1),
	.datab(!cp_ready),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\load_next_out_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam load_next_out_cmd.extended_lut = "off";
defparam load_next_out_cmd.lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam load_next_out_cmd.shared_arith = "off";

dffeas \state.ST_IDLE (
	.clk(clk_clk),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_IDLE~q ),
	.prn(vcc));
defparam \state.ST_IDLE .is_wysiwyg = "true";
defparam \state.ST_IDLE .power_up = "low";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!nxt_out_eop),
	.datac(!stateST_UNCOMP_WR_SUBBURST),
	.datad(!\state.ST_IDLE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'h00EC00EC00EC00EC;
defparam \Selector2~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~1 (
	.dataa(!in_ready_hold),
	.datab(!Equal5),
	.datac(!Equal9),
	.datad(!sink0_data[68]),
	.datae(!src9_valid),
	.dataf(!\Selector2~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~1 .extended_lut = "off";
defparam \Selector2~1 .lut_mask = 64'h0000000100000000;
defparam \Selector2~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~2 (
	.dataa(!\WideOr0~combout ),
	.datab(!\Selector2~1_combout ),
	.datac(!\in_valid~combout ),
	.datad(!nxt_out_eop),
	.datae(!\state.ST_UNCOMP_TRANS~q ),
	.dataf(!sink0_data[69]),
	.datag(!stateST_UNCOMP_WR_SUBBURST),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~2 .extended_lut = "on";
defparam \Selector2~2 .lut_mask = 64'h3B33BB3F0A00AA00;
defparam \Selector2~2 .shared_arith = "off";

dffeas \state.ST_UNCOMP_TRANS (
	.clk(clk_clk),
	.d(\Selector2~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_UNCOMP_TRANS~q ),
	.prn(vcc));
defparam \state.ST_UNCOMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_TRANS .power_up = "low";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!nxt_out_eop),
	.datac(!\state.ST_UNCOMP_TRANS~q ),
	.datad(!stateST_UNCOMP_WR_SUBBURST),
	.datae(!\state.ST_IDLE~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'h0000A8880000A888;
defparam \Selector1~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~1 (
	.dataa(!sink0_data[69]),
	.datab(!stateST_COMP_TRANS),
	.datac(!nxt_out_eop),
	.datad(!sink0_data[68]),
	.datae(!\in_valid~combout ),
	.dataf(!\Selector1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~1 .extended_lut = "off";
defparam \Selector1~1 .lut_mask = 64'h3030777530303330;
defparam \Selector1~1 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[3] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[3]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[3]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[3] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[3] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[2]~2 (
	.dataa(!h2f_ARLEN_0),
	.datab(!sink0_data[69]),
	.datac(!sink0_data[68]),
	.datad(!write_cp_data_74),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[2]~2 .extended_lut = "off";
defparam \d0_int_bytes_remaining[2]~2 .lut_mask = 64'h2F222F222F222F22;
defparam \d0_int_bytes_remaining[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[2]~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\int_bytes_remaining_reg[2]~q ),
	.datad(!\d0_int_bytes_remaining[2]~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[2]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[2]~3 .extended_lut = "off";
defparam \d0_int_bytes_remaining[2]~3 .lut_mask = 64'h287D287D287D287D;
defparam \d0_int_bytes_remaining[2]~3 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[2] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[2]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[2]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[2] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[3]~0 (
	.dataa(!sink0_data[69]),
	.datab(!sink0_data[68]),
	.datac(!write_cp_data_75),
	.datad(!Add2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[3]~0 .extended_lut = "off";
defparam \d0_int_bytes_remaining[3]~0 .lut_mask = 64'h0357035703570357;
defparam \d0_int_bytes_remaining[3]~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[3]~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\int_bytes_remaining_reg[3]~q ),
	.datac(!out_byte_cnt_reg_2),
	.datad(!\int_bytes_remaining_reg[2]~q ),
	.datae(!\d0_int_bytes_remaining[3]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[3]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[3]~1 .extended_lut = "off";
defparam \d0_int_bytes_remaining[3]~1 .lut_mask = 64'h28227D7728227D77;
defparam \d0_int_bytes_remaining[3]~1 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[6] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[6]~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[6]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[6] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[6] .power_up = "low";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!\int_bytes_remaining_reg[3]~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\int_bytes_remaining_reg[2]~q ),
	.datad(!\int_bytes_remaining_reg[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'hDF20DF20DF20DF20;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[4]~8 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!sink0_data[68]),
	.datad(!write_cp_data_76),
	.datae(!Add21),
	.dataf(!\Add1~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[4]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[4]~8 .extended_lut = "off";
defparam \d0_int_bytes_remaining[4]~8 .lut_mask = 64'hCCCFDDDF00031113;
defparam \d0_int_bytes_remaining[4]~8 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[4] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[4]~8_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[4]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[4] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[4] .power_up = "low";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!\int_bytes_remaining_reg[3]~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\int_bytes_remaining_reg[2]~q ),
	.datad(!\int_bytes_remaining_reg[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h2000200020002000;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[5]~6 (
	.dataa(!sink0_data[69]),
	.datab(!sink0_data[68]),
	.datac(!write_cp_data_77),
	.datad(!Add22),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[5]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[5]~6 .extended_lut = "off";
defparam \d0_int_bytes_remaining[5]~6 .lut_mask = 64'h0357035703570357;
defparam \d0_int_bytes_remaining[5]~6 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[5]~7 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\int_bytes_remaining_reg[5]~q ),
	.datac(!\Add1~0_combout ),
	.datad(!\d0_int_bytes_remaining[5]~6_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[5]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[5]~7 .extended_lut = "off";
defparam \d0_int_bytes_remaining[5]~7 .lut_mask = 64'h287D287D287D287D;
defparam \d0_int_bytes_remaining[5]~7 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[5] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[5]~7_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[5]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[5] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[5] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[6]~4 (
	.dataa(!sink0_data[69]),
	.datab(!sink0_data[68]),
	.datac(!write_cp_data_78),
	.datad(!Add23),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[6]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[6]~4 .extended_lut = "off";
defparam \d0_int_bytes_remaining[6]~4 .lut_mask = 64'h0357035703570357;
defparam \d0_int_bytes_remaining[6]~4 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[6]~5 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\int_bytes_remaining_reg[6]~q ),
	.datac(!\int_bytes_remaining_reg[5]~q ),
	.datad(!\Add1~0_combout ),
	.datae(!\d0_int_bytes_remaining[6]~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[6]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[6]~5 .extended_lut = "off";
defparam \d0_int_bytes_remaining[6]~5 .lut_mask = 64'h228277D7228277D7;
defparam \d0_int_bytes_remaining[6]~5 .shared_arith = "off";

cyclonev_lcell_comb \new_burst_reg~0 (
	.dataa(!\Selector1~1_combout ),
	.datab(!\d0_int_bytes_remaining[3]~1_combout ),
	.datac(!\d0_int_bytes_remaining[2]~3_combout ),
	.datad(!\d0_int_bytes_remaining[6]~5_combout ),
	.datae(!\d0_int_bytes_remaining[5]~7_combout ),
	.dataf(!\d0_int_bytes_remaining[4]~8_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\new_burst_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \new_burst_reg~0 .extended_lut = "off";
defparam \new_burst_reg~0 .lut_mask = 64'hAEAAAAAAAAAAAAAA;
defparam \new_burst_reg~0 .shared_arith = "off";

dffeas new_burst_reg(
	.clk(clk_clk),
	.d(\new_burst_reg~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\new_burst_reg~q ),
	.prn(vcc));
defparam new_burst_reg.is_wysiwyg = "true";
defparam new_burst_reg.power_up = "low";

cyclonev_lcell_comb \WideNor0~0 (
	.dataa(!sink0_data[69]),
	.datab(!sink0_data[68]),
	.datac(!WideNor0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideNor0~0 .extended_lut = "off";
defparam \WideNor0~0 .lut_mask = 64'h8A8A8A8A8A8A8A8A;
defparam \WideNor0~0 .shared_arith = "off";

cyclonev_lcell_comb \NON_PIPELINED_INPUTS.load_next_cmd (
	.dataa(!in_ready_hold),
	.datab(!nxt_in_ready1),
	.datac(!nxt_in_ready),
	.datad(!src_valid),
	.datae(!src_valid1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \NON_PIPELINED_INPUTS.load_next_cmd .extended_lut = "off";
defparam \NON_PIPELINED_INPUTS.load_next_cmd .lut_mask = 64'h0015151500151515;
defparam \NON_PIPELINED_INPUTS.load_next_cmd .shared_arith = "off";

dffeas in_bytecount_reg_zero(
	.clk(clk_clk),
	.d(\WideNor0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_bytecount_reg_zero~q ),
	.prn(vcc));
defparam in_bytecount_reg_zero.is_wysiwyg = "true";
defparam in_bytecount_reg_zero.power_up = "low";

cyclonev_lcell_comb \nxt_out_valid~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!\new_burst_reg~q ),
	.datac(!\in_bytecount_reg_zero~q ),
	.datad(!\in_valid~combout ),
	.datae(!cp_ready1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_valid~0 .extended_lut = "off";
defparam \nxt_out_valid~0 .lut_mask = 64'h50FF44FF50FF44FF;
defparam \nxt_out_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!sink0_data[87]),
	.datab(!sink0_data[88]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h8888888888888888;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~0 (
	.dataa(!nxt_out_eop),
	.datab(!\state.ST_UNCOMP_TRANS~q ),
	.datac(!stateST_UNCOMP_WR_SUBBURST),
	.datad(!\WideOr0~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'h002A002A002A002A;
defparam \Selector3~0 .shared_arith = "off";

dffeas \in_size_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[86]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[0]~q ),
	.prn(vcc));
defparam \in_size_reg[0] .is_wysiwyg = "true";
defparam \in_size_reg[0] .power_up = "low";

dffeas \in_size_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[87]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[1]~q ),
	.prn(vcc));
defparam \in_size_reg[1] .is_wysiwyg = "true";
defparam \in_size_reg[1] .power_up = "low";

dffeas \in_size_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[88]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[2]~q ),
	.prn(vcc));
defparam \in_size_reg[2] .is_wysiwyg = "true";
defparam \in_size_reg[2] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[87]),
	.datac(!sink0_data[88]),
	.datad(!\in_size_reg[1]~q ),
	.datae(!\in_size_reg[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~0 .extended_lut = "off";
defparam \ShiftLeft0~0 .lut_mask = 64'h10BA101010BA1010;
defparam \ShiftLeft0~0 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~1 .extended_lut = "off";
defparam \ShiftLeft0~1 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~1 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[3] (
	.clk(clk_clk),
	.d(\ShiftLeft0~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[3]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[3] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[3] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~2 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~2 .extended_lut = "off";
defparam \ShiftLeft0~2 .lut_mask = 64'h00E400E400E400E4;
defparam \ShiftLeft0~2 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[2] (
	.clk(clk_clk),
	.d(\ShiftLeft0~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[2]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[2] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[2] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[87]),
	.datac(!sink0_data[88]),
	.datad(!\in_size_reg[1]~q ),
	.datae(!\in_size_reg[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~3 .extended_lut = "off";
defparam \ShiftLeft0~3 .lut_mask = 64'hEA404040EA404040;
defparam \ShiftLeft0~3 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~4 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~4 .extended_lut = "off";
defparam \ShiftLeft0~4 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~4 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[1] (
	.clk(clk_clk),
	.d(\ShiftLeft0~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[1]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[1] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[1] .power_up = "low";

dffeas \int_byte_cnt_narrow_reg[0] (
	.clk(clk_clk),
	.d(\align_address_to_size|LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[0]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[0] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[0] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[0]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~3 (
	.dataa(!h2f_ARADDR_0),
	.datab(!sink0_data[69]),
	.datac(!sink0_data[68]),
	.datad(!out_data_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~3 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~3 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[0]~3 .shared_arith = "off";

dffeas \in_burstwrap_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[79]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[0]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[0] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[0] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[0]~0 (
	.dataa(!Selector13),
	.datab(!Selector6),
	.datac(!sink0_data[68]),
	.datad(!sink0_data[69]),
	.datae(!\new_burst_reg~q ),
	.dataf(!\d0_int_nxt_addr[0]~4_combout ),
	.datag(!\in_burstwrap_reg[0]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[0]~0 .extended_lut = "on";
defparam \nxt_addr[0]~0 .lut_mask = 64'h00000000F0F0FCA8;
defparam \nxt_addr[0]~0 .shared_arith = "off";

dffeas \int_nxt_addr_reg[0] (
	.clk(clk_clk),
	.d(\nxt_addr[0]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[0] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~4 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\Add0~13_sumout ),
	.datac(!\align_address_to_size|LessThan0~0_combout ),
	.datad(!\d0_int_nxt_addr[0]~3_combout ),
	.datae(!\int_nxt_addr_reg[0]~q ),
	.dataf(!\in_burstwrap_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~4 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~4 .lut_mask = 64'h0005AAAF2227AAAF;
defparam \d0_int_nxt_addr[0]~4 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[0] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[0]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[0] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[1]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[1]~q ),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \in_burstwrap_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[80]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[1]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[1] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[1] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[1]~4 (
	.dataa(!Selector12),
	.datab(!Selector5),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!\new_burst_reg~q ),
	.dataf(!\d0_int_nxt_addr[1]~2_combout ),
	.datag(!\in_burstwrap_reg[1]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[1]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[1]~4 .extended_lut = "on";
defparam \nxt_addr[1]~4 .lut_mask = 64'h00000000F0F0FAC8;
defparam \nxt_addr[1]~4 .shared_arith = "off";

dffeas \int_nxt_addr_reg[1] (
	.clk(clk_clk),
	.d(\nxt_addr[1]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[1] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~7 (
	.dataa(!h2f_ARADDR_1),
	.datab(!sink0_data[69]),
	.datac(!sink0_data[68]),
	.datad(!out_data_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~7 .extended_lut = "off";
defparam \d0_int_nxt_addr[1]~7 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[1]~7 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~2 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\Add0~9_sumout ),
	.datac(!\in_burstwrap_reg[1]~q ),
	.datad(!\int_nxt_addr_reg[1]~q ),
	.datae(!\ShiftLeft0~3_combout ),
	.dataf(!\d0_int_nxt_addr[1]~7_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~2 .extended_lut = "off";
defparam \d0_int_nxt_addr[1]~2 .lut_mask = 64'h02AA02AA02AA57FF;
defparam \d0_int_nxt_addr[1]~2 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[1] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[1]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[1] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_2),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[2]~q ),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[3]~q ),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

dffeas \in_burstwrap_reg[3] (
	.clk(clk_clk),
	.d(sink0_data[82]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[3]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[3] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[3] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[3]~12 (
	.dataa(!Selector10),
	.datab(!Selector3),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!\new_burst_reg~q ),
	.dataf(!\d0_int_nxt_addr[3]~0_combout ),
	.datag(!\in_burstwrap_reg[3]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[3]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[3]~12 .extended_lut = "on";
defparam \nxt_addr[3]~12 .lut_mask = 64'h00000000F0F0FAC8;
defparam \nxt_addr[3]~12 .shared_arith = "off";

dffeas \int_nxt_addr_reg[3] (
	.clk(clk_clk),
	.d(\nxt_addr[3]~12_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[3]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[3] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~5 (
	.dataa(!\Add0~1_sumout ),
	.datab(!\in_burstwrap_reg[3]~q ),
	.datac(!\int_nxt_addr_reg[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~5 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~5 .lut_mask = 64'hE0E0E0E0E0E0E0E0;
defparam \d0_int_nxt_addr[3]~5 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!h2f_ARADDR_3),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!base_address_3),
	.dataf(!\d0_int_nxt_addr[3]~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~0 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~0 .lut_mask = 64'hABABABFF01010155;
defparam \d0_int_nxt_addr[3]~0 .shared_arith = "off";

dffeas \in_burstwrap_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[81]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[2]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[2] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[2] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[2]~8 (
	.dataa(!Selector11),
	.datab(!Selector4),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!\new_burst_reg~q ),
	.dataf(!\d0_int_nxt_addr[2]~1_combout ),
	.datag(!\in_burstwrap_reg[2]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[2]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[2]~8 .extended_lut = "on";
defparam \nxt_addr[2]~8 .lut_mask = 64'h00000000F0F0FAC8;
defparam \nxt_addr[2]~8 .shared_arith = "off";

dffeas \int_nxt_addr_reg[2] (
	.clk(clk_clk),
	.d(\nxt_addr[2]~8_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[2]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~6 (
	.dataa(!\Add0~5_sumout ),
	.datab(!\in_burstwrap_reg[2]~q ),
	.datac(!\int_nxt_addr_reg[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~6 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~6 .lut_mask = 64'hE0E0E0E0E0E0E0E0;
defparam \d0_int_nxt_addr[2]~6 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!h2f_ARADDR_2),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!base_address_2),
	.dataf(!\d0_int_nxt_addr[2]~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~1 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~1 .lut_mask = 64'hABABABFF01010155;
defparam \d0_int_nxt_addr[2]~1 .shared_arith = "off";

dffeas in_eop_reg(
	.clk(clk_clk),
	.d(sink0_endofpacket),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_eop_reg~q ),
	.prn(vcc));
defparam in_eop_reg.is_wysiwyg = "true";
defparam in_eop_reg.power_up = "low";

endmodule

module spw_babasu_altera_merlin_address_alignment_8 (
	new_burst_reg,
	src_data_86,
	in_size_reg_0,
	ShiftLeft0,
	LessThan0)/* synthesis synthesis_greybox=0 */;
input 	new_burst_reg;
input 	src_data_86;
input 	in_size_reg_0;
input 	ShiftLeft0;
output 	LessThan0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!new_burst_reg),
	.datab(!src_data_86),
	.datac(!in_size_reg_0),
	.datad(!ShiftLeft0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan0),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h00E400E400E400E4;
defparam \LessThan0~0 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_burst_adapter_8 (
	h2f_ARADDR_0,
	h2f_ARADDR_1,
	h2f_ARADDR_2,
	h2f_ARADDR_3,
	h2f_ARBURST_0,
	h2f_ARBURST_1,
	h2f_ARID_0,
	h2f_ARID_1,
	h2f_ARID_2,
	h2f_ARID_3,
	h2f_ARID_4,
	h2f_ARID_5,
	h2f_ARID_6,
	h2f_ARID_7,
	h2f_ARID_8,
	h2f_ARID_9,
	h2f_ARID_10,
	h2f_ARID_11,
	h2f_ARLEN_0,
	Add5,
	Add51,
	in_ready_hold,
	saved_grant_1,
	stateST_COMP_TRANS,
	mem_used_1,
	in_data_reg_69,
	in_narrow_reg,
	cp_ready,
	cp_ready1,
	nxt_out_eop,
	out_valid_reg,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready,
	altera_reset_synchronizer_int_chain_out,
	Decoder1,
	Add2,
	Add21,
	Add22,
	Add23,
	src_valid,
	nxt_in_ready1,
	out_byte_cnt_reg_2,
	cp_ready2,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_6,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	Selector10,
	Selector101,
	Selector11,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	Selector12,
	src_payload,
	src_payload1,
	src_payload2,
	Selector13,
	nxt_out_burstwrap_1,
	nxt_addr_2,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARADDR_0;
input 	h2f_ARADDR_1;
input 	h2f_ARADDR_2;
input 	h2f_ARADDR_3;
input 	h2f_ARBURST_0;
input 	h2f_ARBURST_1;
input 	h2f_ARID_0;
input 	h2f_ARID_1;
input 	h2f_ARID_2;
input 	h2f_ARID_3;
input 	h2f_ARID_4;
input 	h2f_ARID_5;
input 	h2f_ARID_6;
input 	h2f_ARID_7;
input 	h2f_ARID_8;
input 	h2f_ARID_9;
input 	h2f_ARID_10;
input 	h2f_ARID_11;
input 	h2f_ARLEN_0;
input 	Add5;
input 	Add51;
input 	in_ready_hold;
input 	saved_grant_1;
output 	stateST_COMP_TRANS;
input 	mem_used_1;
output 	in_data_reg_69;
output 	in_narrow_reg;
input 	cp_ready;
input 	cp_ready1;
output 	nxt_out_eop;
output 	out_valid_reg;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready;
input 	altera_reset_synchronizer_int_chain_out;
input 	Decoder1;
input 	Add2;
input 	Add21;
input 	Add22;
input 	Add23;
input 	src_valid;
output 	nxt_in_ready1;
output 	out_byte_cnt_reg_2;
input 	cp_ready2;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_6;
output 	in_data_reg_105;
output 	in_data_reg_106;
output 	in_data_reg_107;
output 	in_data_reg_108;
output 	in_data_reg_109;
output 	in_data_reg_110;
output 	in_data_reg_111;
output 	in_data_reg_112;
output 	in_data_reg_113;
output 	in_data_reg_114;
output 	in_data_reg_115;
output 	in_data_reg_116;
input 	Selector10;
input 	Selector101;
input 	Selector11;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
input 	Selector12;
input 	src_payload;
input 	src_payload1;
input 	src_payload2;
input 	Selector13;
input 	nxt_out_burstwrap_1;
input 	nxt_addr_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



spw_babasu_altera_merlin_burst_adapter_13_1_8 \altera_merlin_burst_adapter_13_1.burst_adapter (
	.h2f_ARADDR_0(h2f_ARADDR_0),
	.h2f_ARADDR_1(h2f_ARADDR_1),
	.h2f_ARADDR_2(h2f_ARADDR_2),
	.h2f_ARADDR_3(h2f_ARADDR_3),
	.h2f_ARBURST_0(h2f_ARBURST_0),
	.h2f_ARBURST_1(h2f_ARBURST_1),
	.sink0_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,h2f_ARID_11,h2f_ARID_10,h2f_ARID_9,h2f_ARID_8,h2f_ARID_7,h2f_ARID_6,h2f_ARID_5,h2f_ARID_4,h2f_ARID_3,h2f_ARID_2,h2f_ARID_1,h2f_ARID_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_payload2,src_payload1,src_payload,gnd,gnd,gnd,
Selector101,Selector11,Selector12,Selector13,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,saved_grant_1,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.h2f_ARLEN_0(h2f_ARLEN_0),
	.Add5(Add5),
	.Add51(Add51),
	.in_ready_hold(in_ready_hold),
	.stateST_COMP_TRANS(stateST_COMP_TRANS),
	.mem_used_1(mem_used_1),
	.in_data_reg_69(in_data_reg_69),
	.in_narrow_reg1(in_narrow_reg),
	.cp_ready(cp_ready),
	.cp_ready1(cp_ready1),
	.nxt_out_eop(nxt_out_eop),
	.out_valid_reg1(out_valid_reg),
	.stateST_UNCOMP_WR_SUBBURST(stateST_UNCOMP_WR_SUBBURST),
	.nxt_in_ready(nxt_in_ready),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.Decoder1(Decoder1),
	.Add2(Add2),
	.Add21(Add21),
	.Add22(Add22),
	.Add23(Add23),
	.src_valid(src_valid),
	.nxt_in_ready1(nxt_in_ready1),
	.out_byte_cnt_reg_2(out_byte_cnt_reg_2),
	.cp_ready2(cp_ready2),
	.out_uncomp_byte_cnt_reg_5(out_uncomp_byte_cnt_reg_5),
	.out_uncomp_byte_cnt_reg_4(out_uncomp_byte_cnt_reg_4),
	.out_uncomp_byte_cnt_reg_3(out_uncomp_byte_cnt_reg_3),
	.out_uncomp_byte_cnt_reg_2(out_uncomp_byte_cnt_reg_2),
	.out_uncomp_byte_cnt_reg_6(out_uncomp_byte_cnt_reg_6),
	.in_data_reg_105(in_data_reg_105),
	.in_data_reg_106(in_data_reg_106),
	.in_data_reg_107(in_data_reg_107),
	.in_data_reg_108(in_data_reg_108),
	.in_data_reg_109(in_data_reg_109),
	.in_data_reg_110(in_data_reg_110),
	.in_data_reg_111(in_data_reg_111),
	.in_data_reg_112(in_data_reg_112),
	.in_data_reg_113(in_data_reg_113),
	.in_data_reg_114(in_data_reg_114),
	.in_data_reg_115(in_data_reg_115),
	.in_data_reg_116(in_data_reg_116),
	.Selector10(Selector10),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_3),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_2),
	.nxt_out_burstwrap_1(nxt_out_burstwrap_1),
	.nxt_addr_2(nxt_addr_2),
	.clk_clk(clk_clk));

endmodule

module spw_babasu_altera_merlin_burst_adapter_13_1_8 (
	h2f_ARADDR_0,
	h2f_ARADDR_1,
	h2f_ARADDR_2,
	h2f_ARADDR_3,
	h2f_ARBURST_0,
	h2f_ARBURST_1,
	sink0_data,
	h2f_ARLEN_0,
	Add5,
	Add51,
	in_ready_hold,
	stateST_COMP_TRANS,
	mem_used_1,
	in_data_reg_69,
	in_narrow_reg1,
	cp_ready,
	cp_ready1,
	nxt_out_eop,
	out_valid_reg1,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready,
	altera_reset_synchronizer_int_chain_out,
	Decoder1,
	Add2,
	Add21,
	Add22,
	Add23,
	src_valid,
	nxt_in_ready1,
	out_byte_cnt_reg_2,
	cp_ready2,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_6,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	Selector10,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	nxt_out_burstwrap_1,
	nxt_addr_2,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARADDR_0;
input 	h2f_ARADDR_1;
input 	h2f_ARADDR_2;
input 	h2f_ARADDR_3;
input 	h2f_ARBURST_0;
input 	h2f_ARBURST_1;
input 	[128:0] sink0_data;
input 	h2f_ARLEN_0;
input 	Add5;
input 	Add51;
input 	in_ready_hold;
output 	stateST_COMP_TRANS;
input 	mem_used_1;
output 	in_data_reg_69;
output 	in_narrow_reg1;
input 	cp_ready;
input 	cp_ready1;
output 	nxt_out_eop;
output 	out_valid_reg1;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready;
input 	altera_reset_synchronizer_int_chain_out;
input 	Decoder1;
input 	Add2;
input 	Add21;
input 	Add22;
input 	Add23;
input 	src_valid;
output 	nxt_in_ready1;
output 	out_byte_cnt_reg_2;
input 	cp_ready2;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_6;
output 	in_data_reg_105;
output 	in_data_reg_106;
output 	in_data_reg_107;
output 	in_data_reg_108;
output 	in_data_reg_109;
output 	in_data_reg_110;
output 	in_data_reg_111;
output 	in_data_reg_112;
output 	in_data_reg_113;
output 	in_data_reg_114;
output 	in_data_reg_115;
output 	in_data_reg_116;
input 	Selector10;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
input 	nxt_out_burstwrap_1;
input 	nxt_addr_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \align_address_to_size|LessThan0~0_combout ;
wire \align_address_to_size|LessThan0~1_combout ;
wire \nxt_uncomp_subburst_byte_cnt~0_combout ;
wire \Add4~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt[5]~1_combout ;
wire \nxt_uncomp_subburst_byte_cnt[4]~2_combout ;
wire \nxt_uncomp_subburst_byte_cnt[3]~3_combout ;
wire \nxt_uncomp_subburst_byte_cnt[6]~4_combout ;
wire \nxt_uncomp_subburst_byte_cnt[2]~5_combout ;
wire \WideNor1~combout ;
wire \Selector2~1_combout ;
wire \load_next_out_cmd~combout ;
wire \state.ST_UNCOMP_TRANS~q ;
wire \Selector2~0_combout ;
wire \Selector0~0_combout ;
wire \state.ST_IDLE~q ;
wire \Selector1~0_combout ;
wire \Selector1~1_combout ;
wire \NON_PIPELINED_INPUTS.load_next_cmd~0_combout ;
wire \int_bytes_remaining_reg[6]~q ;
wire \d0_int_bytes_remaining[2]~1_combout ;
wire \int_bytes_remaining_reg[2]~q ;
wire \d0_int_bytes_remaining[3]~2_combout ;
wire \int_bytes_remaining_reg[3]~q ;
wire \Add1~1_combout ;
wire \d0_int_bytes_remaining[4]~3_combout ;
wire \int_bytes_remaining_reg[4]~q ;
wire \Add1~0_combout ;
wire \d0_int_bytes_remaining[5]~4_combout ;
wire \int_bytes_remaining_reg[5]~q ;
wire \d0_int_bytes_remaining[6]~0_combout ;
wire \new_burst_reg~0_combout ;
wire \new_burst_reg~q ;
wire \in_bytecount_reg_zero~0_combout ;
wire \in_bytecount_reg_zero~q ;
wire \nxt_out_valid~0_combout ;
wire \nxt_out_valid~1_combout ;
wire \Selector3~0_combout ;
wire \in_burstwrap_reg[3]~q ;
wire \nxt_addr[3]~0_combout ;
wire \nxt_addr[3]~combout ;
wire \int_nxt_addr_reg[3]~q ;
wire \in_size_reg[0]~q ;
wire \in_size_reg[1]~q ;
wire \in_size_reg[2]~q ;
wire \ShiftLeft0~0_combout ;
wire \ShiftLeft0~1_combout ;
wire \int_byte_cnt_narrow_reg[3]~q ;
wire \ShiftLeft0~2_combout ;
wire \int_byte_cnt_narrow_reg[2]~q ;
wire \in_burstwrap_reg[1]~q ;
wire \nxt_addr[1]~combout ;
wire \int_nxt_addr_reg[1]~q ;
wire \ShiftLeft0~3_combout ;
wire \int_byte_cnt_narrow_reg[1]~q ;
wire \int_byte_cnt_narrow_reg[0]~q ;
wire \Add0~13_sumout ;
wire \in_burstwrap_reg[0]~q ;
wire \nxt_addr[0]~combout ;
wire \int_nxt_addr_reg[0]~q ;
wire \d0_int_nxt_addr[0]~2_combout ;
wire \d0_int_nxt_addr[0]~3_combout ;
wire \int_nxt_addr_reg_dly[0]~q ;
wire \Add0~14 ;
wire \Add0~9_sumout ;
wire \d0_int_nxt_addr[1]~4_combout ;
wire \int_nxt_addr_reg_dly[1]~q ;
wire \Add0~10 ;
wire \Add0~6 ;
wire \Add0~1_sumout ;
wire \d0_int_nxt_addr[3]~0_combout ;
wire \in_burstwrap_reg[2]~q ;
wire \nxt_addr[2]~1_combout ;
wire \nxt_addr[2]~combout ;
wire \int_nxt_addr_reg[2]~q ;
wire \Add0~5_sumout ;
wire \d0_int_nxt_addr[2]~1_combout ;


spw_babasu_altera_merlin_address_alignment_9 align_address_to_size(
	.new_burst_reg(\new_burst_reg~q ),
	.src_payload(sink0_data[86]),
	.in_size_reg_0(\in_size_reg[0]~q ),
	.src_payload1(sink0_data[87]),
	.in_size_reg_1(\in_size_reg[1]~q ),
	.src_payload2(sink0_data[88]),
	.in_size_reg_2(\in_size_reg[2]~q ),
	.LessThan0(\align_address_to_size|LessThan0~0_combout ),
	.LessThan01(\align_address_to_size|LessThan0~1_combout ));

dffeas \state.ST_COMP_TRANS (
	.clk(clk_clk),
	.d(\Selector1~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_COMP_TRANS),
	.prn(vcc));
defparam \state.ST_COMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_COMP_TRANS .power_up = "low";

dffeas \in_data_reg[69] (
	.clk(clk_clk),
	.d(sink0_data[69]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_69),
	.prn(vcc));
defparam \in_data_reg[69] .is_wysiwyg = "true";
defparam \in_data_reg[69] .power_up = "low";

dffeas in_narrow_reg(
	.clk(clk_clk),
	.d(Decoder1),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_narrow_reg1),
	.prn(vcc));
defparam in_narrow_reg.is_wysiwyg = "true";
defparam in_narrow_reg.power_up = "low";

cyclonev_lcell_comb \nxt_out_eop~0 (
	.dataa(!in_data_reg_69),
	.datab(!stateST_COMP_TRANS),
	.datac(!\new_burst_reg~q ),
	.datad(!mem_used_1),
	.datae(!cp_ready),
	.dataf(!\in_bytecount_reg_zero~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_out_eop),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_eop~0 .extended_lut = "off";
defparam \nxt_out_eop~0 .lut_mask = 64'h4444474477774777;
defparam \nxt_out_eop~0 .shared_arith = "off";

dffeas out_valid_reg(
	.clk(clk_clk),
	.d(\nxt_out_valid~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_valid_reg1),
	.prn(vcc));
defparam out_valid_reg.is_wysiwyg = "true";
defparam out_valid_reg.power_up = "low";

dffeas \state.ST_UNCOMP_WR_SUBBURST (
	.clk(clk_clk),
	.d(\Selector3~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_UNCOMP_WR_SUBBURST),
	.prn(vcc));
defparam \state.ST_UNCOMP_WR_SUBBURST .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_WR_SUBBURST .power_up = "low";

cyclonev_lcell_comb \nxt_in_ready~0 (
	.dataa(!in_ready_hold),
	.datab(!stateST_COMP_TRANS),
	.datac(!mem_used_1),
	.datad(!cp_ready),
	.datae(!out_valid_reg1),
	.dataf(!\Selector2~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~0 .extended_lut = "off";
defparam \nxt_in_ready~0 .lut_mask = 64'h0000FF3F8888BBBB;
defparam \nxt_in_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_in_ready~1 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!cp_ready1),
	.datac(!nxt_out_eop),
	.datad(!nxt_in_ready),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~1 .extended_lut = "off";
defparam \nxt_in_ready~1 .lut_mask = 64'h00FE00FE00FE00FE;
defparam \nxt_in_ready~1 .shared_arith = "off";

dffeas \out_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[5] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[5]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_5),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[5] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[5] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[4] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[4]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_4),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[4] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[4] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[3] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[3]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_3),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[3] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[3] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[2]~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[6] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[6]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_6),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[6] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[6] .power_up = "low";

dffeas \in_data_reg[105] (
	.clk(clk_clk),
	.d(sink0_data[105]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_105),
	.prn(vcc));
defparam \in_data_reg[105] .is_wysiwyg = "true";
defparam \in_data_reg[105] .power_up = "low";

dffeas \in_data_reg[106] (
	.clk(clk_clk),
	.d(sink0_data[106]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_106),
	.prn(vcc));
defparam \in_data_reg[106] .is_wysiwyg = "true";
defparam \in_data_reg[106] .power_up = "low";

dffeas \in_data_reg[107] (
	.clk(clk_clk),
	.d(sink0_data[107]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_107),
	.prn(vcc));
defparam \in_data_reg[107] .is_wysiwyg = "true";
defparam \in_data_reg[107] .power_up = "low";

dffeas \in_data_reg[108] (
	.clk(clk_clk),
	.d(sink0_data[108]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_108),
	.prn(vcc));
defparam \in_data_reg[108] .is_wysiwyg = "true";
defparam \in_data_reg[108] .power_up = "low";

dffeas \in_data_reg[109] (
	.clk(clk_clk),
	.d(sink0_data[109]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_109),
	.prn(vcc));
defparam \in_data_reg[109] .is_wysiwyg = "true";
defparam \in_data_reg[109] .power_up = "low";

dffeas \in_data_reg[110] (
	.clk(clk_clk),
	.d(sink0_data[110]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_110),
	.prn(vcc));
defparam \in_data_reg[110] .is_wysiwyg = "true";
defparam \in_data_reg[110] .power_up = "low";

dffeas \in_data_reg[111] (
	.clk(clk_clk),
	.d(sink0_data[111]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_111),
	.prn(vcc));
defparam \in_data_reg[111] .is_wysiwyg = "true";
defparam \in_data_reg[111] .power_up = "low";

dffeas \in_data_reg[112] (
	.clk(clk_clk),
	.d(sink0_data[112]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_112),
	.prn(vcc));
defparam \in_data_reg[112] .is_wysiwyg = "true";
defparam \in_data_reg[112] .power_up = "low";

dffeas \in_data_reg[113] (
	.clk(clk_clk),
	.d(sink0_data[113]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_113),
	.prn(vcc));
defparam \in_data_reg[113] .is_wysiwyg = "true";
defparam \in_data_reg[113] .power_up = "low";

dffeas \in_data_reg[114] (
	.clk(clk_clk),
	.d(sink0_data[114]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_114),
	.prn(vcc));
defparam \in_data_reg[114] .is_wysiwyg = "true";
defparam \in_data_reg[114] .power_up = "low";

dffeas \in_data_reg[115] (
	.clk(clk_clk),
	.d(sink0_data[115]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_115),
	.prn(vcc));
defparam \in_data_reg[115] .is_wysiwyg = "true";
defparam \in_data_reg[115] .power_up = "low";

dffeas \in_data_reg[116] (
	.clk(clk_clk),
	.d(sink0_data[116]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_116),
	.prn(vcc));
defparam \in_data_reg[116] .is_wysiwyg = "true";
defparam \in_data_reg[116] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[3] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[3]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_3),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[3] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[2] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[2]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_2),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[2] .power_up = "low";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt~0 (
	.dataa(!cp_ready1),
	.datab(!out_valid_reg1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt~0 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt~0 .lut_mask = 64'h1111111111111111;
defparam \nxt_uncomp_subburst_byte_cnt~0 .shared_arith = "off";

cyclonev_lcell_comb \Add4~0 (
	.dataa(!out_uncomp_byte_cnt_reg_4),
	.datab(!out_uncomp_byte_cnt_reg_3),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add4~0 .extended_lut = "off";
defparam \Add4~0 .lut_mask = 64'h0800080008000800;
defparam \Add4~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[5]~1 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!\Add4~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[5]~1 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[5]~1 .lut_mask = 64'h0F4EA5E40F4EA5E4;
defparam \nxt_uncomp_subburst_byte_cnt[5]~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[4]~2 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!out_uncomp_byte_cnt_reg_3),
	.datae(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.dataf(!out_uncomp_byte_cnt_reg_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[4]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[4]~2 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[4]~2 .lut_mask = 64'h0F0FE44E0F0F4E4E;
defparam \nxt_uncomp_subburst_byte_cnt[4]~2 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[3]~3 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!out_uncomp_byte_cnt_reg_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[3]~3 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[3]~3 .lut_mask = 64'h0FE40F4E0FE40F4E;
defparam \nxt_uncomp_subburst_byte_cnt[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[6]~4 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!\Add4~0_combout ),
	.dataf(!out_uncomp_byte_cnt_reg_6),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[6]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[6]~4 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[6]~4 .lut_mask = 64'h0044A0E4FFEE5F4E;
defparam \nxt_uncomp_subburst_byte_cnt[6]~4 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[2]~5 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[2]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[2]~5 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[2]~5 .lut_mask = 64'h0EF40EF40EF40EF4;
defparam \nxt_uncomp_subburst_byte_cnt[2]~5 .shared_arith = "off";

cyclonev_lcell_comb WideNor1(
	.dataa(!\nxt_uncomp_subburst_byte_cnt[5]~1_combout ),
	.datab(!\nxt_uncomp_subburst_byte_cnt[4]~2_combout ),
	.datac(!\nxt_uncomp_subburst_byte_cnt[3]~3_combout ),
	.datad(!\nxt_uncomp_subburst_byte_cnt[6]~4_combout ),
	.datae(!\nxt_uncomp_subburst_byte_cnt[2]~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideNor1.extended_lut = "off";
defparam WideNor1.lut_mask = 64'h8000000080000000;
defparam WideNor1.shared_arith = "off";

cyclonev_lcell_comb \Selector2~1 (
	.dataa(!nxt_out_eop),
	.datab(!\Selector2~0_combout ),
	.datac(!\WideNor1~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~1 .extended_lut = "off";
defparam \Selector2~1 .lut_mask = 64'h0808080808080808;
defparam \Selector2~1 .shared_arith = "off";

cyclonev_lcell_comb load_next_out_cmd(
	.dataa(!mem_used_1),
	.datab(!cp_ready),
	.datac(!out_valid_reg1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\load_next_out_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam load_next_out_cmd.extended_lut = "off";
defparam load_next_out_cmd.lut_mask = 64'hF2F2F2F2F2F2F2F2;
defparam load_next_out_cmd.shared_arith = "off";

dffeas \state.ST_UNCOMP_TRANS (
	.clk(clk_clk),
	.d(\Selector2~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_UNCOMP_TRANS~q ),
	.prn(vcc));
defparam \state.ST_UNCOMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_TRANS .power_up = "low";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'h8888888888888888;
defparam \Selector2~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!in_ready_hold),
	.datab(!nxt_out_eop),
	.datac(!src_valid),
	.datad(!\state.ST_IDLE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'h05CD05CD05CD05CD;
defparam \Selector0~0 .shared_arith = "off";

dffeas \state.ST_IDLE (
	.clk(clk_clk),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_IDLE~q ),
	.prn(vcc));
defparam \state.ST_IDLE .is_wysiwyg = "true";
defparam \state.ST_IDLE .power_up = "low";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!sink0_data[69]),
	.datab(!nxt_out_eop),
	.datac(!\Selector2~0_combout ),
	.datad(!\state.ST_IDLE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'h5510551055105510;
defparam \Selector1~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~1 (
	.dataa(!in_ready_hold),
	.datab(!stateST_COMP_TRANS),
	.datac(!nxt_out_eop),
	.datad(!src_valid),
	.datae(!\Selector1~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~1 .extended_lut = "off";
defparam \Selector1~1 .lut_mask = 64'h3031307530313075;
defparam \Selector1~1 .shared_arith = "off";

cyclonev_lcell_comb \NON_PIPELINED_INPUTS.load_next_cmd~0 (
	.dataa(!in_ready_hold),
	.datab(!nxt_in_ready1),
	.datac(!src_valid),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \NON_PIPELINED_INPUTS.load_next_cmd~0 .extended_lut = "off";
defparam \NON_PIPELINED_INPUTS.load_next_cmd~0 .lut_mask = 64'h0404040404040404;
defparam \NON_PIPELINED_INPUTS.load_next_cmd~0 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[6] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[6]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[6]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[6] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[6] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[2]~1 (
	.dataa(!h2f_ARLEN_0),
	.datab(!sink0_data[69]),
	.datac(!\new_burst_reg~q ),
	.datad(!out_byte_cnt_reg_2),
	.datae(!\int_bytes_remaining_reg[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[2]~1 .extended_lut = "off";
defparam \d0_int_bytes_remaining[2]~1 .lut_mask = 64'h02F2F20202F2F202;
defparam \d0_int_bytes_remaining[2]~1 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[2] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[2]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[2]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[2] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[3]~2 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!Add2),
	.datad(!\int_bytes_remaining_reg[3]~q ),
	.datae(!out_byte_cnt_reg_2),
	.dataf(!\int_bytes_remaining_reg[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[3]~2 .extended_lut = "off";
defparam \d0_int_bytes_remaining[3]~2 .lut_mask = 64'h01CDCD0101CD01CD;
defparam \d0_int_bytes_remaining[3]~2 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[3] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[3]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[3]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[3] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[3] .power_up = "low";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!\int_bytes_remaining_reg[4]~q ),
	.datab(!\int_bytes_remaining_reg[3]~q ),
	.datac(!out_byte_cnt_reg_2),
	.datad(!\int_bytes_remaining_reg[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'hA6AAA6AAA6AAA6AA;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[4]~3 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!Add21),
	.datad(!\Add1~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[4]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[4]~3 .extended_lut = "off";
defparam \d0_int_bytes_remaining[4]~3 .lut_mask = 64'hCD01CD01CD01CD01;
defparam \d0_int_bytes_remaining[4]~3 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[4] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[4]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[4]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[4] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[4] .power_up = "low";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!\int_bytes_remaining_reg[4]~q ),
	.datab(!\int_bytes_remaining_reg[3]~q ),
	.datac(!out_byte_cnt_reg_2),
	.datad(!\int_bytes_remaining_reg[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h0800080008000800;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[5]~4 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!Add22),
	.datad(!\int_bytes_remaining_reg[5]~q ),
	.datae(!\Add1~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[5]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[5]~4 .extended_lut = "off";
defparam \d0_int_bytes_remaining[5]~4 .lut_mask = 64'h01CDCD0101CDCD01;
defparam \d0_int_bytes_remaining[5]~4 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[5] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[5]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[5]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[5] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[5] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[6]~0 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!Add23),
	.datad(!\int_bytes_remaining_reg[6]~q ),
	.datae(!\int_bytes_remaining_reg[5]~q ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[6]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[6]~0 .extended_lut = "off";
defparam \d0_int_bytes_remaining[6]~0 .lut_mask = 64'h01CD01CDCD0101CD;
defparam \d0_int_bytes_remaining[6]~0 .shared_arith = "off";

cyclonev_lcell_comb \new_burst_reg~0 (
	.dataa(!\Selector1~1_combout ),
	.datab(!\d0_int_bytes_remaining[6]~0_combout ),
	.datac(!\d0_int_bytes_remaining[2]~1_combout ),
	.datad(!\d0_int_bytes_remaining[3]~2_combout ),
	.datae(!\d0_int_bytes_remaining[4]~3_combout ),
	.dataf(!\d0_int_bytes_remaining[5]~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\new_burst_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \new_burst_reg~0 .extended_lut = "off";
defparam \new_burst_reg~0 .lut_mask = 64'hAEAAAAAAAAAAAAAA;
defparam \new_burst_reg~0 .shared_arith = "off";

dffeas new_burst_reg(
	.clk(clk_clk),
	.d(\new_burst_reg~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\new_burst_reg~q ),
	.prn(vcc));
defparam new_burst_reg.is_wysiwyg = "true";
defparam new_burst_reg.power_up = "low";

cyclonev_lcell_comb \in_bytecount_reg_zero~0 (
	.dataa(!sink0_data[69]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\in_bytecount_reg_zero~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \in_bytecount_reg_zero~0 .extended_lut = "off";
defparam \in_bytecount_reg_zero~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \in_bytecount_reg_zero~0 .shared_arith = "off";

dffeas in_bytecount_reg_zero(
	.clk(clk_clk),
	.d(\in_bytecount_reg_zero~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_bytecount_reg_zero~q ),
	.prn(vcc));
defparam in_bytecount_reg_zero.is_wysiwyg = "true";
defparam in_bytecount_reg_zero.power_up = "low";

cyclonev_lcell_comb \nxt_out_valid~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!mem_used_1),
	.datac(!\in_bytecount_reg_zero~q ),
	.datad(!cp_ready2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_valid~0 .extended_lut = "off";
defparam \nxt_out_valid~0 .lut_mask = 64'hF0B8F0B8F0B8F0B8;
defparam \nxt_out_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_out_valid~1 (
	.dataa(!in_ready_hold),
	.datab(!stateST_COMP_TRANS),
	.datac(!src_valid),
	.datad(!\nxt_out_valid~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_valid~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_valid~1 .extended_lut = "off";
defparam \nxt_out_valid~1 .lut_mask = 64'h0537053705370537;
defparam \nxt_out_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~0 (
	.dataa(!nxt_out_eop),
	.datab(!\Selector2~0_combout ),
	.datac(!\WideNor1~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'h8080808080808080;
defparam \Selector3~0 .shared_arith = "off";

dffeas \in_burstwrap_reg[3] (
	.clk(clk_clk),
	.d(sink0_data[82]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_burstwrap_reg[3]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[3] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[3] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[3]~0 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!\in_burstwrap_reg[3]~q ),
	.datad(!\d0_int_nxt_addr[3]~0_combout ),
	.datae(!h2f_ARBURST_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[3]~0 .extended_lut = "off";
defparam \nxt_addr[3]~0 .lut_mask = 64'h00F300E200F300E2;
defparam \nxt_addr[3]~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_addr[3] (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!h2f_ARBURST_1),
	.datad(!Add5),
	.datae(!Selector10),
	.dataf(!\nxt_addr[3]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[3] .extended_lut = "off";
defparam \nxt_addr[3] .lut_mask = 64'h00000000FEEEFFEF;
defparam \nxt_addr[3] .shared_arith = "off";

dffeas \int_nxt_addr_reg[3] (
	.clk(clk_clk),
	.d(\nxt_addr[3]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[3]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[3] .power_up = "low";

dffeas \in_size_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[86]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_size_reg[0]~q ),
	.prn(vcc));
defparam \in_size_reg[0] .is_wysiwyg = "true";
defparam \in_size_reg[0] .power_up = "low";

dffeas \in_size_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[87]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_size_reg[1]~q ),
	.prn(vcc));
defparam \in_size_reg[1] .is_wysiwyg = "true";
defparam \in_size_reg[1] .power_up = "low";

dffeas \in_size_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[88]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_size_reg[2]~q ),
	.prn(vcc));
defparam \in_size_reg[2] .is_wysiwyg = "true";
defparam \in_size_reg[2] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[87]),
	.datac(!\in_size_reg[1]~q ),
	.datad(!sink0_data[88]),
	.datae(!\in_size_reg[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~0 .extended_lut = "off";
defparam \ShiftLeft0~0 .lut_mask = 64'h1B0A11001B0A1100;
defparam \ShiftLeft0~0 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~1 .extended_lut = "off";
defparam \ShiftLeft0~1 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~1 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[3] (
	.clk(clk_clk),
	.d(\ShiftLeft0~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[3]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[3] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[3] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~2 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~2 .extended_lut = "off";
defparam \ShiftLeft0~2 .lut_mask = 64'h00E400E400E400E4;
defparam \ShiftLeft0~2 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[2] (
	.clk(clk_clk),
	.d(\ShiftLeft0~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[2]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[2] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[2] .power_up = "low";

dffeas \in_burstwrap_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[80]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_burstwrap_reg[1]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[1] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[1] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[1] (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!\in_burstwrap_reg[1]~q ),
	.datad(!\d0_int_nxt_addr[1]~4_combout ),
	.datae(!nxt_out_burstwrap_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[1] .extended_lut = "off";
defparam \nxt_addr[1] .lut_mask = 64'h00E200F300E200F3;
defparam \nxt_addr[1] .shared_arith = "off";

dffeas \int_nxt_addr_reg[1] (
	.clk(clk_clk),
	.d(\nxt_addr[1]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[1] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\align_address_to_size|LessThan0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~3 .extended_lut = "off";
defparam \ShiftLeft0~3 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~3 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[1] (
	.clk(clk_clk),
	.d(\ShiftLeft0~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[1]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[1] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[1] .power_up = "low";

dffeas \int_byte_cnt_narrow_reg[0] (
	.clk(clk_clk),
	.d(\align_address_to_size|LessThan0~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[0]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[0] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[0] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[0]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \in_burstwrap_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[79]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_burstwrap_reg[0]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[0] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[0] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[0] (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!sink0_data[79]),
	.datad(!\in_burstwrap_reg[0]~q ),
	.datae(!\d0_int_nxt_addr[0]~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[0] .extended_lut = "off";
defparam \nxt_addr[0] .lut_mask = 64'h0000FE320000FE32;
defparam \nxt_addr[0] .shared_arith = "off";

dffeas \int_nxt_addr_reg[0] (
	.clk(clk_clk),
	.d(\nxt_addr[0]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[0] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~2 (
	.dataa(!\Add0~13_sumout ),
	.datab(!\int_nxt_addr_reg[0]~q ),
	.datac(!\in_burstwrap_reg[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~2 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~2 .lut_mask = 64'hC8C8C8C8C8C8C8C8;
defparam \d0_int_nxt_addr[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~3 (
	.dataa(!h2f_ARADDR_0),
	.datab(!sink0_data[69]),
	.datac(!\new_burst_reg~q ),
	.datad(!\align_address_to_size|LessThan0~1_combout ),
	.datae(!\d0_int_nxt_addr[0]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~3 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~3 .lut_mask = 64'hF0F10001F0F10001;
defparam \d0_int_nxt_addr[0]~3 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[0] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[0]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[0] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[1]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[1]~q ),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~4 (
	.dataa(!\int_nxt_addr_reg[1]~q ),
	.datab(!\Add0~9_sumout ),
	.datac(!sink0_data[69]),
	.datad(!Decoder1),
	.datae(!\new_burst_reg~q ),
	.dataf(!h2f_ARADDR_1),
	.datag(!\in_burstwrap_reg[1]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~4 .extended_lut = "on";
defparam \d0_int_nxt_addr[1]~4 .lut_mask = 64'h575700005757000F;
defparam \d0_int_nxt_addr[1]~4 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[1] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[1]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[1] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_2),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[2]~q ),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[3]~q ),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~0 (
	.dataa(!h2f_ARADDR_3),
	.datab(!sink0_data[69]),
	.datac(!\new_burst_reg~q ),
	.datad(!\int_nxt_addr_reg[3]~q ),
	.datae(!\in_burstwrap_reg[3]~q ),
	.dataf(!\Add0~1_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~0 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~0 .lut_mask = 64'h01F101F101F1F1F1;
defparam \d0_int_nxt_addr[3]~0 .shared_arith = "off";

dffeas \in_burstwrap_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[81]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_burstwrap_reg[2]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[2] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[2] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[2]~1 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!\in_burstwrap_reg[2]~q ),
	.datad(!\d0_int_nxt_addr[2]~1_combout ),
	.datae(!h2f_ARBURST_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[2]~1 .extended_lut = "off";
defparam \nxt_addr[2]~1 .lut_mask = 64'h00F300E200F300E2;
defparam \nxt_addr[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_addr[2] (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!h2f_ARBURST_1),
	.datad(!Add51),
	.datae(!\nxt_addr[2]~1_combout ),
	.dataf(!nxt_addr_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[2] .extended_lut = "off";
defparam \nxt_addr[2] .lut_mask = 64'h0000FEEE0000FFEF;
defparam \nxt_addr[2] .shared_arith = "off";

dffeas \int_nxt_addr_reg[2] (
	.clk(clk_clk),
	.d(\nxt_addr[2]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[2]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~1 (
	.dataa(!h2f_ARADDR_2),
	.datab(!sink0_data[69]),
	.datac(!\new_burst_reg~q ),
	.datad(!\int_nxt_addr_reg[2]~q ),
	.datae(!\in_burstwrap_reg[2]~q ),
	.dataf(!\Add0~5_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~1 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~1 .lut_mask = 64'h01F101F101F1F1F1;
defparam \d0_int_nxt_addr[2]~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_address_alignment_9 (
	new_burst_reg,
	src_payload,
	in_size_reg_0,
	src_payload1,
	in_size_reg_1,
	src_payload2,
	in_size_reg_2,
	LessThan0,
	LessThan01)/* synthesis synthesis_greybox=0 */;
input 	new_burst_reg;
input 	src_payload;
input 	in_size_reg_0;
input 	src_payload1;
input 	in_size_reg_1;
input 	src_payload2;
input 	in_size_reg_2;
output 	LessThan0;
output 	LessThan01;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!new_burst_reg),
	.datab(!src_payload1),
	.datac(!in_size_reg_1),
	.datad(!src_payload2),
	.datae(!in_size_reg_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan0),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'hE4A04400E4A04400;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~1 (
	.dataa(!new_burst_reg),
	.datab(!src_payload),
	.datac(!in_size_reg_0),
	.datad(!LessThan0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan01),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~1 .extended_lut = "off";
defparam \LessThan0~1 .lut_mask = 64'h00E400E400E400E4;
defparam \LessThan0~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_burst_adapter_9 (
	h2f_ARADDR_0,
	h2f_ARADDR_1,
	h2f_ARADDR_2,
	h2f_ARADDR_3,
	h2f_ARLEN_0,
	nxt_in_ready,
	in_ready_hold,
	stateST_COMP_TRANS,
	out_valid_reg,
	mem_used_1,
	in_narrow_reg,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	in_data_reg_68,
	cp_ready,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready1,
	saved_grant_1,
	saved_grant_0,
	altera_reset_synchronizer_int_chain_out,
	in_data_reg_0,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	Add2,
	Add21,
	Add22,
	Add23,
	write_cp_data_77,
	write_cp_data_78,
	write_cp_data_75,
	write_cp_data_74,
	write_cp_data_76,
	WideNor0,
	nxt_out_eop,
	src_valid,
	src_valid1,
	WideOr1,
	cp_ready1,
	cp_ready2,
	in_data_reg_69,
	src_data_87,
	src_data_88,
	src_data_35,
	src_data_34,
	src_data_33,
	src_data_32,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_6,
	src_payload_0,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	Selector3,
	Selector10,
	base_address_3,
	Selector4,
	Selector11,
	base_address_2,
	src_payload,
	src_data_82,
	src_data_81,
	src_data_105,
	src_data_106,
	src_data_107,
	src_data_108,
	src_data_109,
	src_data_110,
	src_data_111,
	src_data_112,
	src_data_113,
	src_data_114,
	src_data_115,
	src_data_116,
	src_data_86,
	Selector5,
	Selector12,
	out_data_1,
	src_data_80,
	out_data_0,
	Selector6,
	Selector13,
	src_data_79,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARADDR_0;
input 	h2f_ARADDR_1;
input 	h2f_ARADDR_2;
input 	h2f_ARADDR_3;
input 	h2f_ARLEN_0;
output 	nxt_in_ready;
input 	in_ready_hold;
output 	stateST_COMP_TRANS;
output 	out_valid_reg;
input 	mem_used_1;
output 	in_narrow_reg;
output 	in_byteen_reg_3;
output 	in_byteen_reg_2;
output 	in_byteen_reg_1;
output 	in_byteen_reg_0;
output 	in_data_reg_68;
input 	cp_ready;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready1;
input 	saved_grant_1;
input 	saved_grant_0;
input 	altera_reset_synchronizer_int_chain_out;
output 	in_data_reg_0;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
input 	Add2;
input 	Add21;
input 	Add22;
input 	Add23;
input 	write_cp_data_77;
input 	write_cp_data_78;
input 	write_cp_data_75;
input 	write_cp_data_74;
input 	write_cp_data_76;
input 	WideNor0;
output 	nxt_out_eop;
input 	src_valid;
input 	src_valid1;
input 	WideOr1;
input 	cp_ready1;
input 	cp_ready2;
output 	in_data_reg_69;
input 	src_data_87;
input 	src_data_88;
input 	src_data_35;
input 	src_data_34;
input 	src_data_33;
input 	src_data_32;
output 	out_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_6;
input 	src_payload_0;
output 	in_data_reg_105;
output 	in_data_reg_106;
output 	in_data_reg_107;
output 	in_data_reg_108;
output 	in_data_reg_109;
output 	in_data_reg_110;
output 	in_data_reg_111;
output 	in_data_reg_112;
output 	in_data_reg_113;
output 	in_data_reg_114;
output 	in_data_reg_115;
output 	in_data_reg_116;
input 	Selector3;
input 	Selector10;
input 	base_address_3;
input 	Selector4;
input 	Selector11;
input 	base_address_2;
input 	src_payload;
input 	src_data_82;
input 	src_data_81;
input 	src_data_105;
input 	src_data_106;
input 	src_data_107;
input 	src_data_108;
input 	src_data_109;
input 	src_data_110;
input 	src_data_111;
input 	src_data_112;
input 	src_data_113;
input 	src_data_114;
input 	src_data_115;
input 	src_data_116;
input 	src_data_86;
input 	Selector5;
input 	Selector12;
input 	out_data_1;
input 	src_data_80;
input 	out_data_0;
input 	Selector6;
input 	Selector13;
input 	src_data_79;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



spw_babasu_altera_merlin_burst_adapter_13_1_9 \altera_merlin_burst_adapter_13_1.burst_adapter (
	.h2f_ARADDR_0(h2f_ARADDR_0),
	.h2f_ARADDR_1(h2f_ARADDR_1),
	.h2f_ARADDR_2(h2f_ARADDR_2),
	.h2f_ARADDR_3(h2f_ARADDR_3),
	.h2f_ARLEN_0(h2f_ARLEN_0),
	.nxt_in_ready(nxt_in_ready),
	.in_ready_hold(in_ready_hold),
	.stateST_COMP_TRANS(stateST_COMP_TRANS),
	.out_valid_reg1(out_valid_reg),
	.mem_used_1(mem_used_1),
	.in_narrow_reg1(in_narrow_reg),
	.in_byteen_reg_3(in_byteen_reg_3),
	.in_byteen_reg_2(in_byteen_reg_2),
	.in_byteen_reg_1(in_byteen_reg_1),
	.in_byteen_reg_0(in_byteen_reg_0),
	.in_data_reg_68(in_data_reg_68),
	.cp_ready(cp_ready),
	.stateST_UNCOMP_WR_SUBBURST(stateST_UNCOMP_WR_SUBBURST),
	.nxt_in_ready1(nxt_in_ready1),
	.sink0_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_116,src_data_115,src_data_114,src_data_113,src_data_112,src_data_111,src_data_110,src_data_109,src_data_108,src_data_107,src_data_106,src_data_105,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_88,src_data_87,
src_data_86,gnd,gnd,gnd,src_data_82,src_data_81,src_data_80,src_data_79,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,saved_grant_1,saved_grant_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_35,src_data_34,src_data_33,
src_data_32,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_payload}),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.in_data_reg_0(in_data_reg_0),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_3),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_2),
	.Add2(Add2),
	.Add21(Add21),
	.Add22(Add22),
	.Add23(Add23),
	.write_cp_data_77(write_cp_data_77),
	.write_cp_data_78(write_cp_data_78),
	.write_cp_data_75(write_cp_data_75),
	.write_cp_data_74(write_cp_data_74),
	.write_cp_data_76(write_cp_data_76),
	.WideNor0(WideNor0),
	.nxt_out_eop(nxt_out_eop),
	.src_valid(src_valid),
	.src_valid1(src_valid1),
	.WideOr1(WideOr1),
	.cp_ready1(cp_ready1),
	.cp_ready2(cp_ready2),
	.in_data_reg_69(in_data_reg_69),
	.out_byte_cnt_reg_2(out_byte_cnt_reg_2),
	.out_uncomp_byte_cnt_reg_5(out_uncomp_byte_cnt_reg_5),
	.out_uncomp_byte_cnt_reg_4(out_uncomp_byte_cnt_reg_4),
	.out_uncomp_byte_cnt_reg_3(out_uncomp_byte_cnt_reg_3),
	.out_uncomp_byte_cnt_reg_2(out_uncomp_byte_cnt_reg_2),
	.out_uncomp_byte_cnt_reg_6(out_uncomp_byte_cnt_reg_6),
	.sink0_endofpacket(src_payload_0),
	.in_data_reg_105(in_data_reg_105),
	.in_data_reg_106(in_data_reg_106),
	.in_data_reg_107(in_data_reg_107),
	.in_data_reg_108(in_data_reg_108),
	.in_data_reg_109(in_data_reg_109),
	.in_data_reg_110(in_data_reg_110),
	.in_data_reg_111(in_data_reg_111),
	.in_data_reg_112(in_data_reg_112),
	.in_data_reg_113(in_data_reg_113),
	.in_data_reg_114(in_data_reg_114),
	.in_data_reg_115(in_data_reg_115),
	.in_data_reg_116(in_data_reg_116),
	.Selector3(Selector3),
	.Selector10(Selector10),
	.base_address_3(base_address_3),
	.Selector4(Selector4),
	.Selector11(Selector11),
	.base_address_2(base_address_2),
	.Selector5(Selector5),
	.Selector12(Selector12),
	.out_data_1(out_data_1),
	.out_data_0(out_data_0),
	.Selector6(Selector6),
	.Selector13(Selector13),
	.clk_clk(clk_clk));

endmodule

module spw_babasu_altera_merlin_burst_adapter_13_1_9 (
	h2f_ARADDR_0,
	h2f_ARADDR_1,
	h2f_ARADDR_2,
	h2f_ARADDR_3,
	h2f_ARLEN_0,
	nxt_in_ready,
	in_ready_hold,
	stateST_COMP_TRANS,
	out_valid_reg1,
	mem_used_1,
	in_narrow_reg1,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	in_data_reg_68,
	cp_ready,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready1,
	sink0_data,
	altera_reset_synchronizer_int_chain_out,
	in_data_reg_0,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	Add2,
	Add21,
	Add22,
	Add23,
	write_cp_data_77,
	write_cp_data_78,
	write_cp_data_75,
	write_cp_data_74,
	write_cp_data_76,
	WideNor0,
	nxt_out_eop,
	src_valid,
	src_valid1,
	WideOr1,
	cp_ready1,
	cp_ready2,
	in_data_reg_69,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_6,
	sink0_endofpacket,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	Selector3,
	Selector10,
	base_address_3,
	Selector4,
	Selector11,
	base_address_2,
	Selector5,
	Selector12,
	out_data_1,
	out_data_0,
	Selector6,
	Selector13,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARADDR_0;
input 	h2f_ARADDR_1;
input 	h2f_ARADDR_2;
input 	h2f_ARADDR_3;
input 	h2f_ARLEN_0;
output 	nxt_in_ready;
input 	in_ready_hold;
output 	stateST_COMP_TRANS;
output 	out_valid_reg1;
input 	mem_used_1;
output 	in_narrow_reg1;
output 	in_byteen_reg_3;
output 	in_byteen_reg_2;
output 	in_byteen_reg_1;
output 	in_byteen_reg_0;
output 	in_data_reg_68;
input 	cp_ready;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready1;
input 	[128:0] sink0_data;
input 	altera_reset_synchronizer_int_chain_out;
output 	in_data_reg_0;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
input 	Add2;
input 	Add21;
input 	Add22;
input 	Add23;
input 	write_cp_data_77;
input 	write_cp_data_78;
input 	write_cp_data_75;
input 	write_cp_data_74;
input 	write_cp_data_76;
input 	WideNor0;
output 	nxt_out_eop;
input 	src_valid;
input 	src_valid1;
input 	WideOr1;
input 	cp_ready1;
input 	cp_ready2;
output 	in_data_reg_69;
output 	out_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_6;
input 	sink0_endofpacket;
output 	in_data_reg_105;
output 	in_data_reg_106;
output 	in_data_reg_107;
output 	in_data_reg_108;
output 	in_data_reg_109;
output 	in_data_reg_110;
output 	in_data_reg_111;
output 	in_data_reg_112;
output 	in_data_reg_113;
output 	in_data_reg_114;
output 	in_data_reg_115;
output 	in_data_reg_116;
input 	Selector3;
input 	Selector10;
input 	base_address_3;
input 	Selector4;
input 	Selector11;
input 	base_address_2;
input 	Selector5;
input 	Selector12;
input 	out_data_1;
input 	out_data_0;
input 	Selector6;
input 	Selector13;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \align_address_to_size|LessThan0~0_combout ;
wire \nxt_in_ready~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt~0_combout ;
wire \Add4~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt[5]~1_combout ;
wire \nxt_uncomp_subburst_byte_cnt[4]~2_combout ;
wire \nxt_uncomp_subburst_byte_cnt[3]~3_combout ;
wire \nxt_uncomp_subburst_byte_cnt[2]~4_combout ;
wire \nxt_uncomp_subburst_byte_cnt[6]~5_combout ;
wire \WideOr0~combout ;
wire \Selector0~0_combout ;
wire \load_next_out_cmd~combout ;
wire \state.ST_IDLE~q ;
wire \Selector2~0_combout ;
wire \Selector2~1_combout ;
wire \Selector2~2_combout ;
wire \state.ST_UNCOMP_TRANS~q ;
wire \Selector1~3_combout ;
wire \Selector1~4_combout ;
wire \Selector1~5_combout ;
wire \int_bytes_remaining_reg[6]~q ;
wire \d0_int_bytes_remaining[2]~5_combout ;
wire \d0_int_bytes_remaining[2]~6_combout ;
wire \int_bytes_remaining_reg[2]~q ;
wire \d0_int_bytes_remaining[3]~7_combout ;
wire \d0_int_bytes_remaining[3]~8_combout ;
wire \int_bytes_remaining_reg[3]~q ;
wire \Add1~1_combout ;
wire \d0_int_bytes_remaining[4]~4_combout ;
wire \int_bytes_remaining_reg[4]~q ;
wire \Add1~0_combout ;
wire \d0_int_bytes_remaining[5]~2_combout ;
wire \d0_int_bytes_remaining[5]~3_combout ;
wire \int_bytes_remaining_reg[5]~q ;
wire \d0_int_bytes_remaining[6]~0_combout ;
wire \d0_int_bytes_remaining[6]~1_combout ;
wire \Equal0~0_combout ;
wire \new_burst_reg~0_combout ;
wire \new_burst_reg~q ;
wire \Selector1~0_combout ;
wire \Selector1~1_combout ;
wire \Selector1~2_combout ;
wire \WideNor0~0_combout ;
wire \NON_PIPELINED_INPUTS.load_next_cmd~combout ;
wire \in_bytecount_reg_zero~q ;
wire \nxt_out_valid~0_combout ;
wire \nxt_out_valid~1_combout ;
wire \LessThan0~0_combout ;
wire \Selector3~0_combout ;
wire \in_size_reg[0]~q ;
wire \in_size_reg[2]~q ;
wire \in_size_reg[1]~q ;
wire \ShiftLeft0~0_combout ;
wire \ShiftLeft0~1_combout ;
wire \int_byte_cnt_narrow_reg[3]~q ;
wire \ShiftLeft0~2_combout ;
wire \int_byte_cnt_narrow_reg[2]~q ;
wire \ShiftLeft0~3_combout ;
wire \ShiftLeft0~4_combout ;
wire \int_byte_cnt_narrow_reg[1]~q ;
wire \int_byte_cnt_narrow_reg[0]~q ;
wire \Add0~13_sumout ;
wire \d0_int_nxt_addr[0]~3_combout ;
wire \in_burstwrap_reg[0]~q ;
wire \nxt_addr[0]~0_combout ;
wire \int_nxt_addr_reg[0]~q ;
wire \d0_int_nxt_addr[0]~4_combout ;
wire \int_nxt_addr_reg_dly[0]~q ;
wire \Add0~14 ;
wire \Add0~9_sumout ;
wire \in_burstwrap_reg[1]~q ;
wire \nxt_addr[1]~4_combout ;
wire \int_nxt_addr_reg[1]~q ;
wire \d0_int_nxt_addr[1]~7_combout ;
wire \d0_int_nxt_addr[1]~2_combout ;
wire \int_nxt_addr_reg_dly[1]~q ;
wire \Add0~10 ;
wire \Add0~6 ;
wire \Add0~1_sumout ;
wire \in_burstwrap_reg[3]~q ;
wire \nxt_addr[3]~12_combout ;
wire \int_nxt_addr_reg[3]~q ;
wire \d0_int_nxt_addr[3]~5_combout ;
wire \d0_int_nxt_addr[3]~0_combout ;
wire \Add0~5_sumout ;
wire \in_burstwrap_reg[2]~q ;
wire \nxt_addr[2]~8_combout ;
wire \int_nxt_addr_reg[2]~q ;
wire \d0_int_nxt_addr[2]~6_combout ;
wire \d0_int_nxt_addr[2]~1_combout ;
wire \in_eop_reg~q ;


spw_babasu_altera_merlin_address_alignment_10 align_address_to_size(
	.new_burst_reg(\new_burst_reg~q ),
	.src_data_86(sink0_data[86]),
	.in_size_reg_0(\in_size_reg[0]~q ),
	.ShiftLeft0(\ShiftLeft0~3_combout ),
	.LessThan0(\align_address_to_size|LessThan0~0_combout ));

cyclonev_lcell_comb \nxt_in_ready~2 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!in_ready_hold),
	.datac(!out_valid_reg1),
	.datad(!cp_ready),
	.datae(!stateST_COMP_TRANS),
	.dataf(!\new_burst_reg~q ),
	.datag(!stateST_UNCOMP_WR_SUBBURST),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~2 .extended_lut = "on";
defparam \nxt_in_ready~2 .lut_mask = 64'h2020F0F02020F0FF;
defparam \nxt_in_ready~2 .shared_arith = "off";

dffeas \state.ST_COMP_TRANS (
	.clk(clk_clk),
	.d(\Selector1~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_COMP_TRANS),
	.prn(vcc));
defparam \state.ST_COMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_COMP_TRANS .power_up = "low";

dffeas out_valid_reg(
	.clk(clk_clk),
	.d(\nxt_out_valid~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_valid_reg1),
	.prn(vcc));
defparam out_valid_reg.is_wysiwyg = "true";
defparam out_valid_reg.power_up = "low";

dffeas in_narrow_reg(
	.clk(clk_clk),
	.d(\LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_narrow_reg1),
	.prn(vcc));
defparam in_narrow_reg.is_wysiwyg = "true";
defparam in_narrow_reg.power_up = "low";

dffeas \in_byteen_reg[3] (
	.clk(clk_clk),
	.d(sink0_data[35]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_3),
	.prn(vcc));
defparam \in_byteen_reg[3] .is_wysiwyg = "true";
defparam \in_byteen_reg[3] .power_up = "low";

dffeas \in_byteen_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[34]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_2),
	.prn(vcc));
defparam \in_byteen_reg[2] .is_wysiwyg = "true";
defparam \in_byteen_reg[2] .power_up = "low";

dffeas \in_byteen_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[33]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_1),
	.prn(vcc));
defparam \in_byteen_reg[1] .is_wysiwyg = "true";
defparam \in_byteen_reg[1] .power_up = "low";

dffeas \in_byteen_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[32]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_0),
	.prn(vcc));
defparam \in_byteen_reg[0] .is_wysiwyg = "true";
defparam \in_byteen_reg[0] .power_up = "low";

dffeas \in_data_reg[68] (
	.clk(clk_clk),
	.d(sink0_data[68]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_68),
	.prn(vcc));
defparam \in_data_reg[68] .is_wysiwyg = "true";
defparam \in_data_reg[68] .power_up = "low";

dffeas \state.ST_UNCOMP_WR_SUBBURST (
	.clk(clk_clk),
	.d(\Selector3~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_UNCOMP_WR_SUBBURST),
	.prn(vcc));
defparam \state.ST_UNCOMP_WR_SUBBURST .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_WR_SUBBURST .power_up = "low";

cyclonev_lcell_comb \nxt_in_ready~1 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!out_valid_reg1),
	.datac(!cp_ready),
	.datad(!\nxt_in_ready~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~1 .extended_lut = "off";
defparam \nxt_in_ready~1 .lut_mask = 64'h8A008A008A008A00;
defparam \nxt_in_ready~1 .shared_arith = "off";

dffeas \in_data_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[0]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_0),
	.prn(vcc));
defparam \in_data_reg[0] .is_wysiwyg = "true";
defparam \in_data_reg[0] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[3] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[3]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_3),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[3] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[2] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[2]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_2),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[2] .power_up = "low";

cyclonev_lcell_comb \nxt_out_eop~0 (
	.dataa(!\in_eop_reg~q ),
	.datab(!stateST_COMP_TRANS),
	.datac(!\new_burst_reg~q ),
	.datad(!cp_ready),
	.datae(!\in_bytecount_reg_zero~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_out_eop),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_eop~0 .extended_lut = "off";
defparam \nxt_out_eop~0 .lut_mask = 64'h4447774744477747;
defparam \nxt_out_eop~0 .shared_arith = "off";

dffeas \in_data_reg[69] (
	.clk(clk_clk),
	.d(sink0_data[69]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_69),
	.prn(vcc));
defparam \in_data_reg[69] .is_wysiwyg = "true";
defparam \in_data_reg[69] .power_up = "low";

dffeas \out_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[5] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[5]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_5),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[5] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[5] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[4] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[4]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_4),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[4] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[4] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[3] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[3]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_3),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[3] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[3] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[2]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[6] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[6]~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_6),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[6] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[6] .power_up = "low";

dffeas \in_data_reg[105] (
	.clk(clk_clk),
	.d(sink0_data[105]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_105),
	.prn(vcc));
defparam \in_data_reg[105] .is_wysiwyg = "true";
defparam \in_data_reg[105] .power_up = "low";

dffeas \in_data_reg[106] (
	.clk(clk_clk),
	.d(sink0_data[106]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_106),
	.prn(vcc));
defparam \in_data_reg[106] .is_wysiwyg = "true";
defparam \in_data_reg[106] .power_up = "low";

dffeas \in_data_reg[107] (
	.clk(clk_clk),
	.d(sink0_data[107]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_107),
	.prn(vcc));
defparam \in_data_reg[107] .is_wysiwyg = "true";
defparam \in_data_reg[107] .power_up = "low";

dffeas \in_data_reg[108] (
	.clk(clk_clk),
	.d(sink0_data[108]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_108),
	.prn(vcc));
defparam \in_data_reg[108] .is_wysiwyg = "true";
defparam \in_data_reg[108] .power_up = "low";

dffeas \in_data_reg[109] (
	.clk(clk_clk),
	.d(sink0_data[109]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_109),
	.prn(vcc));
defparam \in_data_reg[109] .is_wysiwyg = "true";
defparam \in_data_reg[109] .power_up = "low";

dffeas \in_data_reg[110] (
	.clk(clk_clk),
	.d(sink0_data[110]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_110),
	.prn(vcc));
defparam \in_data_reg[110] .is_wysiwyg = "true";
defparam \in_data_reg[110] .power_up = "low";

dffeas \in_data_reg[111] (
	.clk(clk_clk),
	.d(sink0_data[111]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_111),
	.prn(vcc));
defparam \in_data_reg[111] .is_wysiwyg = "true";
defparam \in_data_reg[111] .power_up = "low";

dffeas \in_data_reg[112] (
	.clk(clk_clk),
	.d(sink0_data[112]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_112),
	.prn(vcc));
defparam \in_data_reg[112] .is_wysiwyg = "true";
defparam \in_data_reg[112] .power_up = "low";

dffeas \in_data_reg[113] (
	.clk(clk_clk),
	.d(sink0_data[113]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_113),
	.prn(vcc));
defparam \in_data_reg[113] .is_wysiwyg = "true";
defparam \in_data_reg[113] .power_up = "low";

dffeas \in_data_reg[114] (
	.clk(clk_clk),
	.d(sink0_data[114]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_114),
	.prn(vcc));
defparam \in_data_reg[114] .is_wysiwyg = "true";
defparam \in_data_reg[114] .power_up = "low";

dffeas \in_data_reg[115] (
	.clk(clk_clk),
	.d(sink0_data[115]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_115),
	.prn(vcc));
defparam \in_data_reg[115] .is_wysiwyg = "true";
defparam \in_data_reg[115] .power_up = "low";

dffeas \in_data_reg[116] (
	.clk(clk_clk),
	.d(sink0_data[116]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_116),
	.prn(vcc));
defparam \in_data_reg[116] .is_wysiwyg = "true";
defparam \in_data_reg[116] .power_up = "low";

cyclonev_lcell_comb \nxt_in_ready~0 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_in_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~0 .extended_lut = "off";
defparam \nxt_in_ready~0 .lut_mask = 64'h8888888888888888;
defparam \nxt_in_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt~0 (
	.dataa(!out_valid_reg1),
	.datab(!cp_ready),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt~0 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt~0 .lut_mask = 64'h1111111111111111;
defparam \nxt_uncomp_subburst_byte_cnt~0 .shared_arith = "off";

cyclonev_lcell_comb \Add4~0 (
	.dataa(!out_uncomp_byte_cnt_reg_4),
	.datab(!out_uncomp_byte_cnt_reg_3),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add4~0 .extended_lut = "off";
defparam \Add4~0 .lut_mask = 64'h0800080008000800;
defparam \Add4~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[5]~1 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!\Add4~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[5]~1 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[5]~1 .lut_mask = 64'h0F4EA5E40F4EA5E4;
defparam \nxt_uncomp_subburst_byte_cnt[5]~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[4]~2 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!out_uncomp_byte_cnt_reg_3),
	.datae(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.dataf(!out_uncomp_byte_cnt_reg_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[4]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[4]~2 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[4]~2 .lut_mask = 64'h0F0FE44E0F0F4E4E;
defparam \nxt_uncomp_subburst_byte_cnt[4]~2 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[3]~3 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!out_uncomp_byte_cnt_reg_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[3]~3 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[3]~3 .lut_mask = 64'h0FE40F4E0FE40F4E;
defparam \nxt_uncomp_subburst_byte_cnt[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[2]~4 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[2]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[2]~4 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[2]~4 .lut_mask = 64'h0EF40EF40EF40EF4;
defparam \nxt_uncomp_subburst_byte_cnt[2]~4 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[6]~5 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!\Add4~0_combout ),
	.dataf(!out_uncomp_byte_cnt_reg_6),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[6]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[6]~5 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[6]~5 .lut_mask = 64'h0044A0E4FFEE5F4E;
defparam \nxt_uncomp_subburst_byte_cnt[6]~5 .shared_arith = "off";

cyclonev_lcell_comb WideOr0(
	.dataa(!\nxt_uncomp_subburst_byte_cnt[5]~1_combout ),
	.datab(!\nxt_uncomp_subburst_byte_cnt[4]~2_combout ),
	.datac(!\nxt_uncomp_subburst_byte_cnt[3]~3_combout ),
	.datad(!\nxt_uncomp_subburst_byte_cnt[2]~4_combout ),
	.datae(!\nxt_uncomp_subburst_byte_cnt[6]~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr0.extended_lut = "off";
defparam WideOr0.lut_mask = 64'h8000000080000000;
defparam WideOr0.shared_arith = "off";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!in_ready_hold),
	.datab(!sink0_data[69]),
	.datac(!nxt_out_eop),
	.datad(!sink0_data[68]),
	.datae(!WideOr1),
	.dataf(!\state.ST_IDLE~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'h11550000F5F5F0F0;
defparam \Selector0~0 .shared_arith = "off";

cyclonev_lcell_comb load_next_out_cmd(
	.dataa(!out_valid_reg1),
	.datab(!cp_ready),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\load_next_out_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam load_next_out_cmd.extended_lut = "off";
defparam load_next_out_cmd.lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam load_next_out_cmd.shared_arith = "off";

dffeas \state.ST_IDLE (
	.clk(clk_clk),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_IDLE~q ),
	.prn(vcc));
defparam \state.ST_IDLE .is_wysiwyg = "true";
defparam \state.ST_IDLE .power_up = "low";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!nxt_out_eop),
	.datac(!stateST_UNCOMP_WR_SUBBURST),
	.datad(!\state.ST_IDLE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'h00EC00EC00EC00EC;
defparam \Selector2~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~1 (
	.dataa(!in_ready_hold),
	.datab(!nxt_out_eop),
	.datac(!\state.ST_UNCOMP_TRANS~q ),
	.datad(!src_valid),
	.datae(!src_valid1),
	.dataf(!\Selector2~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~1 .extended_lut = "off";
defparam \Selector2~1 .lut_mask = 64'h0001555500010101;
defparam \Selector2~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~2 (
	.dataa(!sink0_data[69]),
	.datab(!nxt_out_eop),
	.datac(!\nxt_in_ready~0_combout ),
	.datad(!\WideOr0~combout ),
	.datae(!\Selector2~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~2 .extended_lut = "off";
defparam \Selector2~2 .lut_mask = 64'h00C0AAEA00C0AAEA;
defparam \Selector2~2 .shared_arith = "off";

dffeas \state.ST_UNCOMP_TRANS (
	.clk(clk_clk),
	.d(\Selector2~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_UNCOMP_TRANS~q ),
	.prn(vcc));
defparam \state.ST_UNCOMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_TRANS .power_up = "low";

cyclonev_lcell_comb \Selector1~3 (
	.dataa(!in_ready_hold),
	.datab(!stateST_COMP_TRANS),
	.datac(!nxt_out_eop),
	.datad(!sink0_data[68]),
	.datae(gnd),
	.dataf(!src_valid),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~3 .extended_lut = "off";
defparam \Selector1~3 .lut_mask = 64'h3030303031303130;
defparam \Selector1~3 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~4 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!nxt_out_eop),
	.datac(!\nxt_in_ready~0_combout ),
	.datad(!\state.ST_IDLE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~4 .extended_lut = "off";
defparam \Selector1~4 .lut_mask = 64'h008A008A008A008A;
defparam \Selector1~4 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~5 (
	.dataa(!in_ready_hold),
	.datab(!sink0_data[69]),
	.datac(!src_valid),
	.datad(!src_valid1),
	.datae(!\Selector1~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~5 .extended_lut = "off";
defparam \Selector1~5 .lut_mask = 64'h0111000001110000;
defparam \Selector1~5 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[6] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[6]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[6]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[6] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[6] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[2]~5 (
	.dataa(!h2f_ARLEN_0),
	.datab(!sink0_data[69]),
	.datac(!sink0_data[68]),
	.datad(!write_cp_data_74),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[2]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[2]~5 .extended_lut = "off";
defparam \d0_int_bytes_remaining[2]~5 .lut_mask = 64'h2F222F222F222F22;
defparam \d0_int_bytes_remaining[2]~5 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[2]~6 (
	.dataa(!\new_burst_reg~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\int_bytes_remaining_reg[2]~q ),
	.datad(!\d0_int_bytes_remaining[2]~5_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[2]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[2]~6 .extended_lut = "off";
defparam \d0_int_bytes_remaining[2]~6 .lut_mask = 64'h287D287D287D287D;
defparam \d0_int_bytes_remaining[2]~6 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[2] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[2]~6_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[2]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[2] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[3]~7 (
	.dataa(!sink0_data[69]),
	.datab(!sink0_data[68]),
	.datac(!write_cp_data_75),
	.datad(!Add2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[3]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[3]~7 .extended_lut = "off";
defparam \d0_int_bytes_remaining[3]~7 .lut_mask = 64'h0357035703570357;
defparam \d0_int_bytes_remaining[3]~7 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[3]~8 (
	.dataa(!\new_burst_reg~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\int_bytes_remaining_reg[2]~q ),
	.datad(!\int_bytes_remaining_reg[3]~q ),
	.datae(!\d0_int_bytes_remaining[3]~7_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[3]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[3]~8 .extended_lut = "off";
defparam \d0_int_bytes_remaining[3]~8 .lut_mask = 64'h208A75DF208A75DF;
defparam \d0_int_bytes_remaining[3]~8 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[3] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[3]~8_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[3]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[3] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[3] .power_up = "low";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!out_byte_cnt_reg_2),
	.datab(!\int_bytes_remaining_reg[2]~q ),
	.datac(!\int_bytes_remaining_reg[4]~q ),
	.datad(!\int_bytes_remaining_reg[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'hB4F0B4F0B4F0B4F0;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[4]~4 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!sink0_data[68]),
	.datad(!write_cp_data_76),
	.datae(!Add21),
	.dataf(!\Add1~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[4]~4 .extended_lut = "off";
defparam \d0_int_bytes_remaining[4]~4 .lut_mask = 64'hCCCFDDDF00031113;
defparam \d0_int_bytes_remaining[4]~4 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[4] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[4]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[4]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[4] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[4] .power_up = "low";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!out_byte_cnt_reg_2),
	.datab(!\int_bytes_remaining_reg[2]~q ),
	.datac(!\int_bytes_remaining_reg[4]~q ),
	.datad(!\int_bytes_remaining_reg[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h4000400040004000;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[5]~2 (
	.dataa(!sink0_data[69]),
	.datab(!sink0_data[68]),
	.datac(!write_cp_data_77),
	.datad(!Add22),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[5]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[5]~2 .extended_lut = "off";
defparam \d0_int_bytes_remaining[5]~2 .lut_mask = 64'h0357035703570357;
defparam \d0_int_bytes_remaining[5]~2 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[5]~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\int_bytes_remaining_reg[5]~q ),
	.datac(!\Add1~0_combout ),
	.datad(!\d0_int_bytes_remaining[5]~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[5]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[5]~3 .extended_lut = "off";
defparam \d0_int_bytes_remaining[5]~3 .lut_mask = 64'h287D287D287D287D;
defparam \d0_int_bytes_remaining[5]~3 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[5] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[5]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[5]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[5] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[5] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[6]~0 (
	.dataa(!sink0_data[69]),
	.datab(!sink0_data[68]),
	.datac(!write_cp_data_78),
	.datad(!Add23),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[6]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[6]~0 .extended_lut = "off";
defparam \d0_int_bytes_remaining[6]~0 .lut_mask = 64'h0357035703570357;
defparam \d0_int_bytes_remaining[6]~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[6]~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\int_bytes_remaining_reg[6]~q ),
	.datac(!\int_bytes_remaining_reg[5]~q ),
	.datad(!\Add1~0_combout ),
	.datae(!\d0_int_bytes_remaining[6]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[6]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[6]~1 .extended_lut = "off";
defparam \d0_int_bytes_remaining[6]~1 .lut_mask = 64'h228277D7228277D7;
defparam \d0_int_bytes_remaining[6]~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!\d0_int_bytes_remaining[2]~6_combout ),
	.datab(!\d0_int_bytes_remaining[3]~8_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'h4444444444444444;
defparam \Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \new_burst_reg~0 (
	.dataa(!\Selector1~3_combout ),
	.datab(!\Selector1~5_combout ),
	.datac(!\d0_int_bytes_remaining[6]~1_combout ),
	.datad(!\d0_int_bytes_remaining[5]~3_combout ),
	.datae(!\d0_int_bytes_remaining[4]~4_combout ),
	.dataf(!\Equal0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\new_burst_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \new_burst_reg~0 .extended_lut = "off";
defparam \new_burst_reg~0 .lut_mask = 64'h88888888F8888888;
defparam \new_burst_reg~0 .shared_arith = "off";

dffeas new_burst_reg(
	.clk(clk_clk),
	.d(\new_burst_reg~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\new_burst_reg~q ),
	.prn(vcc));
defparam new_burst_reg.is_wysiwyg = "true";
defparam new_burst_reg.power_up = "low";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!in_ready_hold),
	.datab(!sink0_data[68]),
	.datac(gnd),
	.datad(!src_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'h0044004400440044;
defparam \Selector1~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~1 (
	.dataa(!in_ready_hold),
	.datab(!sink0_data[69]),
	.datac(!src_valid),
	.datad(!src_valid1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~1 .extended_lut = "off";
defparam \Selector1~1 .lut_mask = 64'h0111011101110111;
defparam \Selector1~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~2 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!nxt_out_eop),
	.datac(!\nxt_in_ready~0_combout ),
	.datad(!\state.ST_IDLE~q ),
	.datae(!\Selector1~0_combout ),
	.dataf(!\Selector1~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~2 .extended_lut = "off";
defparam \Selector1~2 .lut_mask = 64'h44445555FF75FF75;
defparam \Selector1~2 .shared_arith = "off";

cyclonev_lcell_comb \WideNor0~0 (
	.dataa(!sink0_data[69]),
	.datab(!sink0_data[68]),
	.datac(!WideNor0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideNor0~0 .extended_lut = "off";
defparam \WideNor0~0 .lut_mask = 64'h8A8A8A8A8A8A8A8A;
defparam \WideNor0~0 .shared_arith = "off";

cyclonev_lcell_comb \NON_PIPELINED_INPUTS.load_next_cmd (
	.dataa(!in_ready_hold),
	.datab(!nxt_in_ready1),
	.datac(!nxt_in_ready),
	.datad(!src_valid),
	.datae(!src_valid1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \NON_PIPELINED_INPUTS.load_next_cmd .extended_lut = "off";
defparam \NON_PIPELINED_INPUTS.load_next_cmd .lut_mask = 64'h0015151500151515;
defparam \NON_PIPELINED_INPUTS.load_next_cmd .shared_arith = "off";

dffeas in_bytecount_reg_zero(
	.clk(clk_clk),
	.d(\WideNor0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_bytecount_reg_zero~q ),
	.prn(vcc));
defparam in_bytecount_reg_zero.is_wysiwyg = "true";
defparam in_bytecount_reg_zero.power_up = "low";

cyclonev_lcell_comb \nxt_out_valid~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!mem_used_1),
	.datac(!\in_bytecount_reg_zero~q ),
	.datad(!cp_ready1),
	.datae(!cp_ready2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_valid~0 .extended_lut = "off";
defparam \nxt_out_valid~0 .lut_mask = 64'hF0B8B8B8F0B8B8B8;
defparam \nxt_out_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_out_valid~1 (
	.dataa(!in_ready_hold),
	.datab(!stateST_COMP_TRANS),
	.datac(!WideOr1),
	.datad(!\nxt_out_valid~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_valid~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_valid~1 .extended_lut = "off";
defparam \nxt_out_valid~1 .lut_mask = 64'h5073507350735073;
defparam \nxt_out_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!sink0_data[87]),
	.datab(!sink0_data[88]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h8888888888888888;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~0 (
	.dataa(!nxt_out_eop),
	.datab(!\nxt_in_ready~0_combout ),
	.datac(!\WideOr0~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'h8080808080808080;
defparam \Selector3~0 .shared_arith = "off";

dffeas \in_size_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[86]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[0]~q ),
	.prn(vcc));
defparam \in_size_reg[0] .is_wysiwyg = "true";
defparam \in_size_reg[0] .power_up = "low";

dffeas \in_size_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[88]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[2]~q ),
	.prn(vcc));
defparam \in_size_reg[2] .is_wysiwyg = "true";
defparam \in_size_reg[2] .power_up = "low";

dffeas \in_size_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[87]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[1]~q ),
	.prn(vcc));
defparam \in_size_reg[1] .is_wysiwyg = "true";
defparam \in_size_reg[1] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[87]),
	.datac(!sink0_data[88]),
	.datad(!\in_size_reg[2]~q ),
	.datae(!\in_size_reg[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~0 .extended_lut = "off";
defparam \ShiftLeft0~0 .lut_mask = 64'h1010BA101010BA10;
defparam \ShiftLeft0~0 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~1 .extended_lut = "off";
defparam \ShiftLeft0~1 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~1 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[3] (
	.clk(clk_clk),
	.d(\ShiftLeft0~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[3]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[3] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[3] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~2 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~2 .extended_lut = "off";
defparam \ShiftLeft0~2 .lut_mask = 64'h00E400E400E400E4;
defparam \ShiftLeft0~2 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[2] (
	.clk(clk_clk),
	.d(\ShiftLeft0~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[2]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[2] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[2] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[87]),
	.datac(!sink0_data[88]),
	.datad(!\in_size_reg[2]~q ),
	.datae(!\in_size_reg[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~3 .extended_lut = "off";
defparam \ShiftLeft0~3 .lut_mask = 64'hEA404040EA404040;
defparam \ShiftLeft0~3 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~4 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~4 .extended_lut = "off";
defparam \ShiftLeft0~4 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~4 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[1] (
	.clk(clk_clk),
	.d(\ShiftLeft0~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[1]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[1] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[1] .power_up = "low";

dffeas \int_byte_cnt_narrow_reg[0] (
	.clk(clk_clk),
	.d(\align_address_to_size|LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[0]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[0] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[0] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[0]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~3 (
	.dataa(!h2f_ARADDR_0),
	.datab(!sink0_data[69]),
	.datac(!sink0_data[68]),
	.datad(!out_data_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~3 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~3 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[0]~3 .shared_arith = "off";

dffeas \in_burstwrap_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[79]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[0]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[0] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[0] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[0]~0 (
	.dataa(!Selector13),
	.datab(!Selector6),
	.datac(!sink0_data[68]),
	.datad(!sink0_data[69]),
	.datae(!\new_burst_reg~q ),
	.dataf(!\d0_int_nxt_addr[0]~4_combout ),
	.datag(!\in_burstwrap_reg[0]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[0]~0 .extended_lut = "on";
defparam \nxt_addr[0]~0 .lut_mask = 64'h00000000F0F0FCA8;
defparam \nxt_addr[0]~0 .shared_arith = "off";

dffeas \int_nxt_addr_reg[0] (
	.clk(clk_clk),
	.d(\nxt_addr[0]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[0] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~4 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\Add0~13_sumout ),
	.datac(!\align_address_to_size|LessThan0~0_combout ),
	.datad(!\d0_int_nxt_addr[0]~3_combout ),
	.datae(!\int_nxt_addr_reg[0]~q ),
	.dataf(!\in_burstwrap_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~4 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~4 .lut_mask = 64'h0005AAAF2227AAAF;
defparam \d0_int_nxt_addr[0]~4 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[0] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[0]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[0] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[1]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[1]~q ),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \in_burstwrap_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[80]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[1]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[1] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[1] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[1]~4 (
	.dataa(!Selector12),
	.datab(!Selector5),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!\new_burst_reg~q ),
	.dataf(!\d0_int_nxt_addr[1]~2_combout ),
	.datag(!\in_burstwrap_reg[1]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[1]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[1]~4 .extended_lut = "on";
defparam \nxt_addr[1]~4 .lut_mask = 64'h00000000F0F0FAC8;
defparam \nxt_addr[1]~4 .shared_arith = "off";

dffeas \int_nxt_addr_reg[1] (
	.clk(clk_clk),
	.d(\nxt_addr[1]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[1] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~7 (
	.dataa(!h2f_ARADDR_1),
	.datab(!sink0_data[69]),
	.datac(!sink0_data[68]),
	.datad(!out_data_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~7 .extended_lut = "off";
defparam \d0_int_nxt_addr[1]~7 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[1]~7 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~2 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\Add0~9_sumout ),
	.datac(!\in_burstwrap_reg[1]~q ),
	.datad(!\int_nxt_addr_reg[1]~q ),
	.datae(!\ShiftLeft0~3_combout ),
	.dataf(!\d0_int_nxt_addr[1]~7_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~2 .extended_lut = "off";
defparam \d0_int_nxt_addr[1]~2 .lut_mask = 64'h02AA02AA02AA57FF;
defparam \d0_int_nxt_addr[1]~2 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[1] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[1]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[1] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_2),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[2]~q ),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[3]~q ),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

dffeas \in_burstwrap_reg[3] (
	.clk(clk_clk),
	.d(sink0_data[82]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[3]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[3] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[3] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[3]~12 (
	.dataa(!Selector10),
	.datab(!Selector3),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!\new_burst_reg~q ),
	.dataf(!\d0_int_nxt_addr[3]~0_combout ),
	.datag(!\in_burstwrap_reg[3]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[3]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[3]~12 .extended_lut = "on";
defparam \nxt_addr[3]~12 .lut_mask = 64'h00000000F0F0FAC8;
defparam \nxt_addr[3]~12 .shared_arith = "off";

dffeas \int_nxt_addr_reg[3] (
	.clk(clk_clk),
	.d(\nxt_addr[3]~12_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[3]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[3] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~5 (
	.dataa(!\Add0~1_sumout ),
	.datab(!\in_burstwrap_reg[3]~q ),
	.datac(!\int_nxt_addr_reg[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~5 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~5 .lut_mask = 64'hE0E0E0E0E0E0E0E0;
defparam \d0_int_nxt_addr[3]~5 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!h2f_ARADDR_3),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!base_address_3),
	.dataf(!\d0_int_nxt_addr[3]~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~0 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~0 .lut_mask = 64'hABABABFF01010155;
defparam \d0_int_nxt_addr[3]~0 .shared_arith = "off";

dffeas \in_burstwrap_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[81]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[2]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[2] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[2] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[2]~8 (
	.dataa(!Selector11),
	.datab(!Selector4),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!\new_burst_reg~q ),
	.dataf(!\d0_int_nxt_addr[2]~1_combout ),
	.datag(!\in_burstwrap_reg[2]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[2]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[2]~8 .extended_lut = "on";
defparam \nxt_addr[2]~8 .lut_mask = 64'h00000000F0F0FAC8;
defparam \nxt_addr[2]~8 .shared_arith = "off";

dffeas \int_nxt_addr_reg[2] (
	.clk(clk_clk),
	.d(\nxt_addr[2]~8_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[2]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~6 (
	.dataa(!\Add0~5_sumout ),
	.datab(!\in_burstwrap_reg[2]~q ),
	.datac(!\int_nxt_addr_reg[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~6 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~6 .lut_mask = 64'hE0E0E0E0E0E0E0E0;
defparam \d0_int_nxt_addr[2]~6 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!h2f_ARADDR_2),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!base_address_2),
	.dataf(!\d0_int_nxt_addr[2]~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~1 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~1 .lut_mask = 64'hABABABFF01010155;
defparam \d0_int_nxt_addr[2]~1 .shared_arith = "off";

dffeas in_eop_reg(
	.clk(clk_clk),
	.d(sink0_endofpacket),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_eop_reg~q ),
	.prn(vcc));
defparam in_eop_reg.is_wysiwyg = "true";
defparam in_eop_reg.power_up = "low";

endmodule

module spw_babasu_altera_merlin_address_alignment_10 (
	new_burst_reg,
	src_data_86,
	in_size_reg_0,
	ShiftLeft0,
	LessThan0)/* synthesis synthesis_greybox=0 */;
input 	new_burst_reg;
input 	src_data_86;
input 	in_size_reg_0;
input 	ShiftLeft0;
output 	LessThan0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!new_burst_reg),
	.datab(!src_data_86),
	.datac(!in_size_reg_0),
	.datad(!ShiftLeft0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan0),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h00E400E400E400E4;
defparam \LessThan0~0 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_burst_adapter_10 (
	h2f_ARADDR_0,
	h2f_ARADDR_1,
	h2f_ARADDR_2,
	h2f_ARADDR_3,
	h2f_ARLEN_0,
	nxt_in_ready,
	in_ready_hold,
	stateST_COMP_TRANS,
	out_valid_reg,
	in_narrow_reg,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	in_data_reg_68,
	cp_ready,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready1,
	saved_grant_1,
	Equal13,
	saved_grant_0,
	altera_reset_synchronizer_int_chain_out,
	in_data_reg_0,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	Add2,
	Add21,
	Add22,
	Add23,
	Equal5,
	write_cp_data_77,
	write_cp_data_78,
	write_cp_data_75,
	write_cp_data_74,
	write_cp_data_76,
	WideNor0,
	nxt_out_eop,
	src13_valid,
	src_valid,
	cp_ready1,
	in_data_reg_69,
	src_data_87,
	src_data_88,
	src_valid1,
	src_data_35,
	src_data_34,
	src_data_33,
	src_data_32,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_6,
	src_payload_0,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	Selector3,
	Selector10,
	base_address_3,
	Selector4,
	Selector11,
	base_address_2,
	src_payload,
	src_data_82,
	src_data_81,
	src_data_105,
	src_data_106,
	src_data_107,
	src_data_108,
	src_data_109,
	src_data_110,
	src_data_111,
	src_data_112,
	src_data_113,
	src_data_114,
	src_data_115,
	src_data_116,
	src_data_86,
	Selector5,
	Selector12,
	out_data_1,
	src_data_80,
	out_data_0,
	Selector6,
	Selector13,
	src_data_79,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARADDR_0;
input 	h2f_ARADDR_1;
input 	h2f_ARADDR_2;
input 	h2f_ARADDR_3;
input 	h2f_ARLEN_0;
output 	nxt_in_ready;
input 	in_ready_hold;
output 	stateST_COMP_TRANS;
output 	out_valid_reg;
output 	in_narrow_reg;
output 	in_byteen_reg_3;
output 	in_byteen_reg_2;
output 	in_byteen_reg_1;
output 	in_byteen_reg_0;
output 	in_data_reg_68;
input 	cp_ready;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready1;
input 	saved_grant_1;
input 	Equal13;
input 	saved_grant_0;
input 	altera_reset_synchronizer_int_chain_out;
output 	in_data_reg_0;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
input 	Add2;
input 	Add21;
input 	Add22;
input 	Add23;
input 	Equal5;
input 	write_cp_data_77;
input 	write_cp_data_78;
input 	write_cp_data_75;
input 	write_cp_data_74;
input 	write_cp_data_76;
input 	WideNor0;
output 	nxt_out_eop;
input 	src13_valid;
input 	src_valid;
input 	cp_ready1;
output 	in_data_reg_69;
input 	src_data_87;
input 	src_data_88;
input 	src_valid1;
input 	src_data_35;
input 	src_data_34;
input 	src_data_33;
input 	src_data_32;
output 	out_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_6;
input 	src_payload_0;
output 	in_data_reg_105;
output 	in_data_reg_106;
output 	in_data_reg_107;
output 	in_data_reg_108;
output 	in_data_reg_109;
output 	in_data_reg_110;
output 	in_data_reg_111;
output 	in_data_reg_112;
output 	in_data_reg_113;
output 	in_data_reg_114;
output 	in_data_reg_115;
output 	in_data_reg_116;
input 	Selector3;
input 	Selector10;
input 	base_address_3;
input 	Selector4;
input 	Selector11;
input 	base_address_2;
input 	src_payload;
input 	src_data_82;
input 	src_data_81;
input 	src_data_105;
input 	src_data_106;
input 	src_data_107;
input 	src_data_108;
input 	src_data_109;
input 	src_data_110;
input 	src_data_111;
input 	src_data_112;
input 	src_data_113;
input 	src_data_114;
input 	src_data_115;
input 	src_data_116;
input 	src_data_86;
input 	Selector5;
input 	Selector12;
input 	out_data_1;
input 	src_data_80;
input 	out_data_0;
input 	Selector6;
input 	Selector13;
input 	src_data_79;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



spw_babasu_altera_merlin_burst_adapter_13_1_10 \altera_merlin_burst_adapter_13_1.burst_adapter (
	.h2f_ARADDR_0(h2f_ARADDR_0),
	.h2f_ARADDR_1(h2f_ARADDR_1),
	.h2f_ARADDR_2(h2f_ARADDR_2),
	.h2f_ARADDR_3(h2f_ARADDR_3),
	.h2f_ARLEN_0(h2f_ARLEN_0),
	.nxt_in_ready(nxt_in_ready),
	.in_ready_hold(in_ready_hold),
	.stateST_COMP_TRANS(stateST_COMP_TRANS),
	.out_valid_reg1(out_valid_reg),
	.in_narrow_reg1(in_narrow_reg),
	.in_byteen_reg_3(in_byteen_reg_3),
	.in_byteen_reg_2(in_byteen_reg_2),
	.in_byteen_reg_1(in_byteen_reg_1),
	.in_byteen_reg_0(in_byteen_reg_0),
	.in_data_reg_68(in_data_reg_68),
	.cp_ready(cp_ready),
	.stateST_UNCOMP_WR_SUBBURST(stateST_UNCOMP_WR_SUBBURST),
	.nxt_in_ready1(nxt_in_ready1),
	.sink0_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_116,src_data_115,src_data_114,src_data_113,src_data_112,src_data_111,src_data_110,src_data_109,src_data_108,src_data_107,src_data_106,src_data_105,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_88,src_data_87,
src_data_86,gnd,gnd,gnd,src_data_82,src_data_81,src_data_80,src_data_79,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,saved_grant_1,saved_grant_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_35,src_data_34,src_data_33,
src_data_32,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_payload}),
	.Equal13(Equal13),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.in_data_reg_0(in_data_reg_0),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_3),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_2),
	.Add2(Add2),
	.Add21(Add21),
	.Add22(Add22),
	.Add23(Add23),
	.Equal5(Equal5),
	.write_cp_data_77(write_cp_data_77),
	.write_cp_data_78(write_cp_data_78),
	.write_cp_data_75(write_cp_data_75),
	.write_cp_data_74(write_cp_data_74),
	.write_cp_data_76(write_cp_data_76),
	.WideNor0(WideNor0),
	.nxt_out_eop(nxt_out_eop),
	.src13_valid(src13_valid),
	.src_valid(src_valid),
	.cp_ready1(cp_ready1),
	.in_data_reg_69(in_data_reg_69),
	.src_valid1(src_valid1),
	.out_byte_cnt_reg_2(out_byte_cnt_reg_2),
	.out_uncomp_byte_cnt_reg_5(out_uncomp_byte_cnt_reg_5),
	.out_uncomp_byte_cnt_reg_4(out_uncomp_byte_cnt_reg_4),
	.out_uncomp_byte_cnt_reg_3(out_uncomp_byte_cnt_reg_3),
	.out_uncomp_byte_cnt_reg_2(out_uncomp_byte_cnt_reg_2),
	.out_uncomp_byte_cnt_reg_6(out_uncomp_byte_cnt_reg_6),
	.sink0_endofpacket(src_payload_0),
	.in_data_reg_105(in_data_reg_105),
	.in_data_reg_106(in_data_reg_106),
	.in_data_reg_107(in_data_reg_107),
	.in_data_reg_108(in_data_reg_108),
	.in_data_reg_109(in_data_reg_109),
	.in_data_reg_110(in_data_reg_110),
	.in_data_reg_111(in_data_reg_111),
	.in_data_reg_112(in_data_reg_112),
	.in_data_reg_113(in_data_reg_113),
	.in_data_reg_114(in_data_reg_114),
	.in_data_reg_115(in_data_reg_115),
	.in_data_reg_116(in_data_reg_116),
	.Selector3(Selector3),
	.Selector10(Selector10),
	.base_address_3(base_address_3),
	.Selector4(Selector4),
	.Selector11(Selector11),
	.base_address_2(base_address_2),
	.Selector5(Selector5),
	.Selector12(Selector12),
	.out_data_1(out_data_1),
	.out_data_0(out_data_0),
	.Selector6(Selector6),
	.Selector13(Selector13),
	.clk_clk(clk_clk));

endmodule

module spw_babasu_altera_merlin_burst_adapter_13_1_10 (
	h2f_ARADDR_0,
	h2f_ARADDR_1,
	h2f_ARADDR_2,
	h2f_ARADDR_3,
	h2f_ARLEN_0,
	nxt_in_ready,
	in_ready_hold,
	stateST_COMP_TRANS,
	out_valid_reg1,
	in_narrow_reg1,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	in_data_reg_68,
	cp_ready,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready1,
	sink0_data,
	Equal13,
	altera_reset_synchronizer_int_chain_out,
	in_data_reg_0,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	Add2,
	Add21,
	Add22,
	Add23,
	Equal5,
	write_cp_data_77,
	write_cp_data_78,
	write_cp_data_75,
	write_cp_data_74,
	write_cp_data_76,
	WideNor0,
	nxt_out_eop,
	src13_valid,
	src_valid,
	cp_ready1,
	in_data_reg_69,
	src_valid1,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_6,
	sink0_endofpacket,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	Selector3,
	Selector10,
	base_address_3,
	Selector4,
	Selector11,
	base_address_2,
	Selector5,
	Selector12,
	out_data_1,
	out_data_0,
	Selector6,
	Selector13,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARADDR_0;
input 	h2f_ARADDR_1;
input 	h2f_ARADDR_2;
input 	h2f_ARADDR_3;
input 	h2f_ARLEN_0;
output 	nxt_in_ready;
input 	in_ready_hold;
output 	stateST_COMP_TRANS;
output 	out_valid_reg1;
output 	in_narrow_reg1;
output 	in_byteen_reg_3;
output 	in_byteen_reg_2;
output 	in_byteen_reg_1;
output 	in_byteen_reg_0;
output 	in_data_reg_68;
input 	cp_ready;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready1;
input 	[128:0] sink0_data;
input 	Equal13;
input 	altera_reset_synchronizer_int_chain_out;
output 	in_data_reg_0;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
input 	Add2;
input 	Add21;
input 	Add22;
input 	Add23;
input 	Equal5;
input 	write_cp_data_77;
input 	write_cp_data_78;
input 	write_cp_data_75;
input 	write_cp_data_74;
input 	write_cp_data_76;
input 	WideNor0;
output 	nxt_out_eop;
input 	src13_valid;
input 	src_valid;
input 	cp_ready1;
output 	in_data_reg_69;
input 	src_valid1;
output 	out_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_6;
input 	sink0_endofpacket;
output 	in_data_reg_105;
output 	in_data_reg_106;
output 	in_data_reg_107;
output 	in_data_reg_108;
output 	in_data_reg_109;
output 	in_data_reg_110;
output 	in_data_reg_111;
output 	in_data_reg_112;
output 	in_data_reg_113;
output 	in_data_reg_114;
output 	in_data_reg_115;
output 	in_data_reg_116;
input 	Selector3;
input 	Selector10;
input 	base_address_3;
input 	Selector4;
input 	Selector11;
input 	base_address_2;
input 	Selector5;
input 	Selector12;
input 	out_data_1;
input 	out_data_0;
input 	Selector6;
input 	Selector13;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \align_address_to_size|LessThan0~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt~0_combout ;
wire \Add4~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt[5]~1_combout ;
wire \nxt_uncomp_subburst_byte_cnt[4]~2_combout ;
wire \nxt_uncomp_subburst_byte_cnt[3]~3_combout ;
wire \nxt_uncomp_subburst_byte_cnt[2]~4_combout ;
wire \nxt_uncomp_subburst_byte_cnt[6]~5_combout ;
wire \WideOr0~combout ;
wire \in_valid~combout ;
wire \Selector0~0_combout ;
wire \load_next_out_cmd~combout ;
wire \state.ST_IDLE~q ;
wire \Selector2~0_combout ;
wire \Selector2~1_combout ;
wire \Selector2~2_combout ;
wire \state.ST_UNCOMP_TRANS~q ;
wire \Selector1~0_combout ;
wire \Selector1~1_combout ;
wire \int_bytes_remaining_reg[5]~q ;
wire \d0_int_bytes_remaining[2]~5_combout ;
wire \d0_int_bytes_remaining[2]~6_combout ;
wire \int_bytes_remaining_reg[2]~q ;
wire \d0_int_bytes_remaining[3]~3_combout ;
wire \d0_int_bytes_remaining[3]~4_combout ;
wire \int_bytes_remaining_reg[3]~q ;
wire \Add1~1_combout ;
wire \d0_int_bytes_remaining[4]~2_combout ;
wire \int_bytes_remaining_reg[4]~q ;
wire \Add1~0_combout ;
wire \d0_int_bytes_remaining[5]~0_combout ;
wire \d0_int_bytes_remaining[5]~1_combout ;
wire \int_bytes_remaining_reg[6]~q ;
wire \d0_int_bytes_remaining[6]~7_combout ;
wire \d0_int_bytes_remaining[6]~8_combout ;
wire \new_burst_reg~0_combout ;
wire \new_burst_reg~q ;
wire \WideNor0~0_combout ;
wire \NON_PIPELINED_INPUTS.load_next_cmd~combout ;
wire \in_bytecount_reg_zero~q ;
wire \nxt_out_valid~0_combout ;
wire \LessThan0~0_combout ;
wire \Selector3~0_combout ;
wire \in_size_reg[0]~q ;
wire \in_size_reg[1]~q ;
wire \in_size_reg[2]~q ;
wire \ShiftLeft0~0_combout ;
wire \ShiftLeft0~1_combout ;
wire \int_byte_cnt_narrow_reg[3]~q ;
wire \ShiftLeft0~2_combout ;
wire \int_byte_cnt_narrow_reg[2]~q ;
wire \ShiftLeft0~3_combout ;
wire \ShiftLeft0~4_combout ;
wire \int_byte_cnt_narrow_reg[1]~q ;
wire \int_byte_cnt_narrow_reg[0]~q ;
wire \Add0~13_sumout ;
wire \d0_int_nxt_addr[0]~3_combout ;
wire \in_burstwrap_reg[0]~q ;
wire \nxt_addr[0]~0_combout ;
wire \int_nxt_addr_reg[0]~q ;
wire \d0_int_nxt_addr[0]~4_combout ;
wire \int_nxt_addr_reg_dly[0]~q ;
wire \Add0~14 ;
wire \Add0~9_sumout ;
wire \in_burstwrap_reg[1]~q ;
wire \nxt_addr[1]~4_combout ;
wire \int_nxt_addr_reg[1]~q ;
wire \d0_int_nxt_addr[1]~7_combout ;
wire \d0_int_nxt_addr[1]~2_combout ;
wire \int_nxt_addr_reg_dly[1]~q ;
wire \Add0~10 ;
wire \Add0~6 ;
wire \Add0~1_sumout ;
wire \in_burstwrap_reg[3]~q ;
wire \nxt_addr[3]~12_combout ;
wire \int_nxt_addr_reg[3]~q ;
wire \d0_int_nxt_addr[3]~5_combout ;
wire \d0_int_nxt_addr[3]~0_combout ;
wire \Add0~5_sumout ;
wire \in_burstwrap_reg[2]~q ;
wire \nxt_addr[2]~8_combout ;
wire \int_nxt_addr_reg[2]~q ;
wire \d0_int_nxt_addr[2]~6_combout ;
wire \d0_int_nxt_addr[2]~1_combout ;
wire \in_eop_reg~q ;


spw_babasu_altera_merlin_address_alignment_11 align_address_to_size(
	.new_burst_reg(\new_burst_reg~q ),
	.src_data_86(sink0_data[86]),
	.in_size_reg_0(\in_size_reg[0]~q ),
	.ShiftLeft0(\ShiftLeft0~3_combout ),
	.LessThan0(\align_address_to_size|LessThan0~0_combout ));

cyclonev_lcell_comb \nxt_in_ready~1 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!in_ready_hold),
	.datac(!out_valid_reg1),
	.datad(!cp_ready),
	.datae(!stateST_COMP_TRANS),
	.dataf(!\new_burst_reg~q ),
	.datag(!stateST_UNCOMP_WR_SUBBURST),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~1 .extended_lut = "on";
defparam \nxt_in_ready~1 .lut_mask = 64'h2020F0F02020F0FF;
defparam \nxt_in_ready~1 .shared_arith = "off";

dffeas \state.ST_COMP_TRANS (
	.clk(clk_clk),
	.d(\Selector1~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_COMP_TRANS),
	.prn(vcc));
defparam \state.ST_COMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_COMP_TRANS .power_up = "low";

dffeas out_valid_reg(
	.clk(clk_clk),
	.d(\nxt_out_valid~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_valid_reg1),
	.prn(vcc));
defparam out_valid_reg.is_wysiwyg = "true";
defparam out_valid_reg.power_up = "low";

dffeas in_narrow_reg(
	.clk(clk_clk),
	.d(\LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_narrow_reg1),
	.prn(vcc));
defparam in_narrow_reg.is_wysiwyg = "true";
defparam in_narrow_reg.power_up = "low";

dffeas \in_byteen_reg[3] (
	.clk(clk_clk),
	.d(sink0_data[35]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_3),
	.prn(vcc));
defparam \in_byteen_reg[3] .is_wysiwyg = "true";
defparam \in_byteen_reg[3] .power_up = "low";

dffeas \in_byteen_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[34]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_2),
	.prn(vcc));
defparam \in_byteen_reg[2] .is_wysiwyg = "true";
defparam \in_byteen_reg[2] .power_up = "low";

dffeas \in_byteen_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[33]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_1),
	.prn(vcc));
defparam \in_byteen_reg[1] .is_wysiwyg = "true";
defparam \in_byteen_reg[1] .power_up = "low";

dffeas \in_byteen_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[32]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_0),
	.prn(vcc));
defparam \in_byteen_reg[0] .is_wysiwyg = "true";
defparam \in_byteen_reg[0] .power_up = "low";

dffeas \in_data_reg[68] (
	.clk(clk_clk),
	.d(sink0_data[68]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_68),
	.prn(vcc));
defparam \in_data_reg[68] .is_wysiwyg = "true";
defparam \in_data_reg[68] .power_up = "low";

dffeas \state.ST_UNCOMP_WR_SUBBURST (
	.clk(clk_clk),
	.d(\Selector3~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_UNCOMP_WR_SUBBURST),
	.prn(vcc));
defparam \state.ST_UNCOMP_WR_SUBBURST .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_WR_SUBBURST .power_up = "low";

cyclonev_lcell_comb \nxt_in_ready~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!out_valid_reg1),
	.datac(!cp_ready),
	.datad(!\state.ST_UNCOMP_TRANS~q ),
	.datae(!stateST_UNCOMP_WR_SUBBURST),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~0 .extended_lut = "off";
defparam \nxt_in_ready~0 .lut_mask = 64'h008A8A8A008A8A8A;
defparam \nxt_in_ready~0 .shared_arith = "off";

dffeas \in_data_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[0]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_0),
	.prn(vcc));
defparam \in_data_reg[0] .is_wysiwyg = "true";
defparam \in_data_reg[0] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[3] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[3]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_3),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[3] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[2] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[2]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_2),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[2] .power_up = "low";

cyclonev_lcell_comb \nxt_out_eop~0 (
	.dataa(!\in_eop_reg~q ),
	.datab(!stateST_COMP_TRANS),
	.datac(!\new_burst_reg~q ),
	.datad(!cp_ready),
	.datae(!\in_bytecount_reg_zero~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_out_eop),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_eop~0 .extended_lut = "off";
defparam \nxt_out_eop~0 .lut_mask = 64'h4447774744477747;
defparam \nxt_out_eop~0 .shared_arith = "off";

dffeas \in_data_reg[69] (
	.clk(clk_clk),
	.d(sink0_data[69]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_69),
	.prn(vcc));
defparam \in_data_reg[69] .is_wysiwyg = "true";
defparam \in_data_reg[69] .power_up = "low";

dffeas \out_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[5] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[5]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_5),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[5] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[5] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[4] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[4]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_4),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[4] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[4] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[3] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[3]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_3),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[3] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[3] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[2]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[6] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[6]~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_6),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[6] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[6] .power_up = "low";

dffeas \in_data_reg[105] (
	.clk(clk_clk),
	.d(sink0_data[105]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_105),
	.prn(vcc));
defparam \in_data_reg[105] .is_wysiwyg = "true";
defparam \in_data_reg[105] .power_up = "low";

dffeas \in_data_reg[106] (
	.clk(clk_clk),
	.d(sink0_data[106]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_106),
	.prn(vcc));
defparam \in_data_reg[106] .is_wysiwyg = "true";
defparam \in_data_reg[106] .power_up = "low";

dffeas \in_data_reg[107] (
	.clk(clk_clk),
	.d(sink0_data[107]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_107),
	.prn(vcc));
defparam \in_data_reg[107] .is_wysiwyg = "true";
defparam \in_data_reg[107] .power_up = "low";

dffeas \in_data_reg[108] (
	.clk(clk_clk),
	.d(sink0_data[108]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_108),
	.prn(vcc));
defparam \in_data_reg[108] .is_wysiwyg = "true";
defparam \in_data_reg[108] .power_up = "low";

dffeas \in_data_reg[109] (
	.clk(clk_clk),
	.d(sink0_data[109]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_109),
	.prn(vcc));
defparam \in_data_reg[109] .is_wysiwyg = "true";
defparam \in_data_reg[109] .power_up = "low";

dffeas \in_data_reg[110] (
	.clk(clk_clk),
	.d(sink0_data[110]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_110),
	.prn(vcc));
defparam \in_data_reg[110] .is_wysiwyg = "true";
defparam \in_data_reg[110] .power_up = "low";

dffeas \in_data_reg[111] (
	.clk(clk_clk),
	.d(sink0_data[111]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_111),
	.prn(vcc));
defparam \in_data_reg[111] .is_wysiwyg = "true";
defparam \in_data_reg[111] .power_up = "low";

dffeas \in_data_reg[112] (
	.clk(clk_clk),
	.d(sink0_data[112]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_112),
	.prn(vcc));
defparam \in_data_reg[112] .is_wysiwyg = "true";
defparam \in_data_reg[112] .power_up = "low";

dffeas \in_data_reg[113] (
	.clk(clk_clk),
	.d(sink0_data[113]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_113),
	.prn(vcc));
defparam \in_data_reg[113] .is_wysiwyg = "true";
defparam \in_data_reg[113] .power_up = "low";

dffeas \in_data_reg[114] (
	.clk(clk_clk),
	.d(sink0_data[114]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_114),
	.prn(vcc));
defparam \in_data_reg[114] .is_wysiwyg = "true";
defparam \in_data_reg[114] .power_up = "low";

dffeas \in_data_reg[115] (
	.clk(clk_clk),
	.d(sink0_data[115]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_115),
	.prn(vcc));
defparam \in_data_reg[115] .is_wysiwyg = "true";
defparam \in_data_reg[115] .power_up = "low";

dffeas \in_data_reg[116] (
	.clk(clk_clk),
	.d(sink0_data[116]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_116),
	.prn(vcc));
defparam \in_data_reg[116] .is_wysiwyg = "true";
defparam \in_data_reg[116] .power_up = "low";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt~0 (
	.dataa(!out_valid_reg1),
	.datab(!cp_ready),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt~0 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt~0 .lut_mask = 64'h1111111111111111;
defparam \nxt_uncomp_subburst_byte_cnt~0 .shared_arith = "off";

cyclonev_lcell_comb \Add4~0 (
	.dataa(!out_uncomp_byte_cnt_reg_4),
	.datab(!out_uncomp_byte_cnt_reg_3),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add4~0 .extended_lut = "off";
defparam \Add4~0 .lut_mask = 64'h0800080008000800;
defparam \Add4~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[5]~1 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!\Add4~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[5]~1 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[5]~1 .lut_mask = 64'h0F4EA5E40F4EA5E4;
defparam \nxt_uncomp_subburst_byte_cnt[5]~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[4]~2 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!out_uncomp_byte_cnt_reg_3),
	.datae(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.dataf(!out_uncomp_byte_cnt_reg_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[4]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[4]~2 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[4]~2 .lut_mask = 64'h0F0FE44E0F0F4E4E;
defparam \nxt_uncomp_subburst_byte_cnt[4]~2 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[3]~3 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!out_uncomp_byte_cnt_reg_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[3]~3 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[3]~3 .lut_mask = 64'h0FE40F4E0FE40F4E;
defparam \nxt_uncomp_subburst_byte_cnt[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[2]~4 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[2]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[2]~4 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[2]~4 .lut_mask = 64'h0EF40EF40EF40EF4;
defparam \nxt_uncomp_subburst_byte_cnt[2]~4 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[6]~5 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!\Add4~0_combout ),
	.dataf(!out_uncomp_byte_cnt_reg_6),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[6]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[6]~5 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[6]~5 .lut_mask = 64'h0044A0E4FFEE5F4E;
defparam \nxt_uncomp_subburst_byte_cnt[6]~5 .shared_arith = "off";

cyclonev_lcell_comb WideOr0(
	.dataa(!\nxt_uncomp_subburst_byte_cnt[5]~1_combout ),
	.datab(!\nxt_uncomp_subburst_byte_cnt[4]~2_combout ),
	.datac(!\nxt_uncomp_subburst_byte_cnt[3]~3_combout ),
	.datad(!\nxt_uncomp_subburst_byte_cnt[2]~4_combout ),
	.datae(!\nxt_uncomp_subburst_byte_cnt[6]~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr0.extended_lut = "off";
defparam WideOr0.lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam WideOr0.shared_arith = "off";

cyclonev_lcell_comb in_valid(
	.dataa(!in_ready_hold),
	.datab(!Equal5),
	.datac(!Equal13),
	.datad(!sink0_data[68]),
	.datae(!src13_valid),
	.dataf(!src_valid),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\in_valid~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam in_valid.extended_lut = "off";
defparam in_valid.lut_mask = 64'h0000000155555555;
defparam in_valid.shared_arith = "off";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!sink0_data[69]),
	.datab(!nxt_out_eop),
	.datac(!sink0_data[68]),
	.datad(!\in_valid~combout ),
	.datae(!\state.ST_IDLE~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'h005FCCFF005FCCFF;
defparam \Selector0~0 .shared_arith = "off";

cyclonev_lcell_comb load_next_out_cmd(
	.dataa(!out_valid_reg1),
	.datab(!cp_ready),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\load_next_out_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam load_next_out_cmd.extended_lut = "off";
defparam load_next_out_cmd.lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam load_next_out_cmd.shared_arith = "off";

dffeas \state.ST_IDLE (
	.clk(clk_clk),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_IDLE~q ),
	.prn(vcc));
defparam \state.ST_IDLE .is_wysiwyg = "true";
defparam \state.ST_IDLE .power_up = "low";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!nxt_out_eop),
	.datac(!stateST_UNCOMP_WR_SUBBURST),
	.datad(!\state.ST_IDLE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'h00EC00EC00EC00EC;
defparam \Selector2~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~1 (
	.dataa(!in_ready_hold),
	.datab(!Equal5),
	.datac(!Equal13),
	.datad(!sink0_data[68]),
	.datae(!src13_valid),
	.dataf(!\Selector2~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~1 .extended_lut = "off";
defparam \Selector2~1 .lut_mask = 64'h0000000100000000;
defparam \Selector2~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~2 (
	.dataa(!\WideOr0~combout ),
	.datab(!\Selector2~1_combout ),
	.datac(!\in_valid~combout ),
	.datad(!nxt_out_eop),
	.datae(!\state.ST_UNCOMP_TRANS~q ),
	.dataf(!sink0_data[69]),
	.datag(!stateST_UNCOMP_WR_SUBBURST),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~2 .extended_lut = "on";
defparam \Selector2~2 .lut_mask = 64'h3B33BB3F0A00AA00;
defparam \Selector2~2 .shared_arith = "off";

dffeas \state.ST_UNCOMP_TRANS (
	.clk(clk_clk),
	.d(\Selector2~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_UNCOMP_TRANS~q ),
	.prn(vcc));
defparam \state.ST_UNCOMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_TRANS .power_up = "low";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!nxt_out_eop),
	.datac(!\state.ST_UNCOMP_TRANS~q ),
	.datad(!stateST_UNCOMP_WR_SUBBURST),
	.datae(!\state.ST_IDLE~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'h0000A8880000A888;
defparam \Selector1~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~1 (
	.dataa(!sink0_data[69]),
	.datab(!stateST_COMP_TRANS),
	.datac(!nxt_out_eop),
	.datad(!sink0_data[68]),
	.datae(!\in_valid~combout ),
	.dataf(!\Selector1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~1 .extended_lut = "off";
defparam \Selector1~1 .lut_mask = 64'h3030777530303330;
defparam \Selector1~1 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[5] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[5]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[5]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[5] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[5] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[2]~5 (
	.dataa(!h2f_ARLEN_0),
	.datab(!sink0_data[69]),
	.datac(!sink0_data[68]),
	.datad(!write_cp_data_74),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[2]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[2]~5 .extended_lut = "off";
defparam \d0_int_bytes_remaining[2]~5 .lut_mask = 64'h2F222F222F222F22;
defparam \d0_int_bytes_remaining[2]~5 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[2]~6 (
	.dataa(!\new_burst_reg~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\int_bytes_remaining_reg[2]~q ),
	.datad(!\d0_int_bytes_remaining[2]~5_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[2]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[2]~6 .extended_lut = "off";
defparam \d0_int_bytes_remaining[2]~6 .lut_mask = 64'h287D287D287D287D;
defparam \d0_int_bytes_remaining[2]~6 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[2] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[2]~6_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[2]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[2] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[3]~3 (
	.dataa(!sink0_data[69]),
	.datab(!sink0_data[68]),
	.datac(!write_cp_data_75),
	.datad(!Add2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[3]~3 .extended_lut = "off";
defparam \d0_int_bytes_remaining[3]~3 .lut_mask = 64'h0357035703570357;
defparam \d0_int_bytes_remaining[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[3]~4 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\int_bytes_remaining_reg[3]~q ),
	.datac(!out_byte_cnt_reg_2),
	.datad(!\int_bytes_remaining_reg[2]~q ),
	.datae(!\d0_int_bytes_remaining[3]~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[3]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[3]~4 .extended_lut = "off";
defparam \d0_int_bytes_remaining[3]~4 .lut_mask = 64'h28227D7728227D77;
defparam \d0_int_bytes_remaining[3]~4 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[3] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[3]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[3]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[3] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[3] .power_up = "low";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!\int_bytes_remaining_reg[4]~q ),
	.datab(!\int_bytes_remaining_reg[3]~q ),
	.datac(!out_byte_cnt_reg_2),
	.datad(!\int_bytes_remaining_reg[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'hA6AAA6AAA6AAA6AA;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[4]~2 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!sink0_data[68]),
	.datad(!write_cp_data_76),
	.datae(!Add21),
	.dataf(!\Add1~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[4]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[4]~2 .extended_lut = "off";
defparam \d0_int_bytes_remaining[4]~2 .lut_mask = 64'hCCCFDDDF00031113;
defparam \d0_int_bytes_remaining[4]~2 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[4] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[4]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[4]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[4] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[4] .power_up = "low";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!\int_bytes_remaining_reg[4]~q ),
	.datab(!\int_bytes_remaining_reg[3]~q ),
	.datac(!out_byte_cnt_reg_2),
	.datad(!\int_bytes_remaining_reg[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h0800080008000800;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[5]~0 (
	.dataa(!sink0_data[69]),
	.datab(!sink0_data[68]),
	.datac(!write_cp_data_77),
	.datad(!Add22),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[5]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[5]~0 .extended_lut = "off";
defparam \d0_int_bytes_remaining[5]~0 .lut_mask = 64'h0357035703570357;
defparam \d0_int_bytes_remaining[5]~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[5]~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\int_bytes_remaining_reg[5]~q ),
	.datac(!\Add1~0_combout ),
	.datad(!\d0_int_bytes_remaining[5]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[5]~1 .extended_lut = "off";
defparam \d0_int_bytes_remaining[5]~1 .lut_mask = 64'h287D287D287D287D;
defparam \d0_int_bytes_remaining[5]~1 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[6] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[6]~8_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[6]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[6] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[6] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[6]~7 (
	.dataa(!sink0_data[69]),
	.datab(!sink0_data[68]),
	.datac(!write_cp_data_78),
	.datad(!Add23),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[6]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[6]~7 .extended_lut = "off";
defparam \d0_int_bytes_remaining[6]~7 .lut_mask = 64'h0357035703570357;
defparam \d0_int_bytes_remaining[6]~7 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[6]~8 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\int_bytes_remaining_reg[5]~q ),
	.datac(!\Add1~0_combout ),
	.datad(!\int_bytes_remaining_reg[6]~q ),
	.datae(!\d0_int_bytes_remaining[6]~7_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[6]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[6]~8 .extended_lut = "off";
defparam \d0_int_bytes_remaining[6]~8 .lut_mask = 64'h08A25DF708A25DF7;
defparam \d0_int_bytes_remaining[6]~8 .shared_arith = "off";

cyclonev_lcell_comb \new_burst_reg~0 (
	.dataa(!\Selector1~1_combout ),
	.datab(!\d0_int_bytes_remaining[5]~1_combout ),
	.datac(!\d0_int_bytes_remaining[4]~2_combout ),
	.datad(!\d0_int_bytes_remaining[3]~4_combout ),
	.datae(!\d0_int_bytes_remaining[2]~6_combout ),
	.dataf(!\d0_int_bytes_remaining[6]~8_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\new_burst_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \new_burst_reg~0 .extended_lut = "off";
defparam \new_burst_reg~0 .lut_mask = 64'hAAAAEAAAAAAAAAAA;
defparam \new_burst_reg~0 .shared_arith = "off";

dffeas new_burst_reg(
	.clk(clk_clk),
	.d(\new_burst_reg~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\new_burst_reg~q ),
	.prn(vcc));
defparam new_burst_reg.is_wysiwyg = "true";
defparam new_burst_reg.power_up = "low";

cyclonev_lcell_comb \WideNor0~0 (
	.dataa(!sink0_data[69]),
	.datab(!sink0_data[68]),
	.datac(!WideNor0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideNor0~0 .extended_lut = "off";
defparam \WideNor0~0 .lut_mask = 64'h8A8A8A8A8A8A8A8A;
defparam \WideNor0~0 .shared_arith = "off";

cyclonev_lcell_comb \NON_PIPELINED_INPUTS.load_next_cmd (
	.dataa(!in_ready_hold),
	.datab(!nxt_in_ready1),
	.datac(!nxt_in_ready),
	.datad(!src_valid),
	.datae(!src_valid1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \NON_PIPELINED_INPUTS.load_next_cmd .extended_lut = "off";
defparam \NON_PIPELINED_INPUTS.load_next_cmd .lut_mask = 64'h0015151500151515;
defparam \NON_PIPELINED_INPUTS.load_next_cmd .shared_arith = "off";

dffeas in_bytecount_reg_zero(
	.clk(clk_clk),
	.d(\WideNor0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_bytecount_reg_zero~q ),
	.prn(vcc));
defparam in_bytecount_reg_zero.is_wysiwyg = "true";
defparam in_bytecount_reg_zero.power_up = "low";

cyclonev_lcell_comb \nxt_out_valid~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!\new_burst_reg~q ),
	.datac(!\in_bytecount_reg_zero~q ),
	.datad(!\in_valid~combout ),
	.datae(!cp_ready1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_valid~0 .extended_lut = "off";
defparam \nxt_out_valid~0 .lut_mask = 64'h50FF44FF50FF44FF;
defparam \nxt_out_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!sink0_data[87]),
	.datab(!sink0_data[88]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h8888888888888888;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~0 (
	.dataa(!nxt_out_eop),
	.datab(!\state.ST_UNCOMP_TRANS~q ),
	.datac(!stateST_UNCOMP_WR_SUBBURST),
	.datad(!\WideOr0~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'h002A002A002A002A;
defparam \Selector3~0 .shared_arith = "off";

dffeas \in_size_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[86]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[0]~q ),
	.prn(vcc));
defparam \in_size_reg[0] .is_wysiwyg = "true";
defparam \in_size_reg[0] .power_up = "low";

dffeas \in_size_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[87]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[1]~q ),
	.prn(vcc));
defparam \in_size_reg[1] .is_wysiwyg = "true";
defparam \in_size_reg[1] .power_up = "low";

dffeas \in_size_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[88]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[2]~q ),
	.prn(vcc));
defparam \in_size_reg[2] .is_wysiwyg = "true";
defparam \in_size_reg[2] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[87]),
	.datac(!sink0_data[88]),
	.datad(!\in_size_reg[1]~q ),
	.datae(!\in_size_reg[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~0 .extended_lut = "off";
defparam \ShiftLeft0~0 .lut_mask = 64'h10BA101010BA1010;
defparam \ShiftLeft0~0 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~1 .extended_lut = "off";
defparam \ShiftLeft0~1 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~1 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[3] (
	.clk(clk_clk),
	.d(\ShiftLeft0~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[3]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[3] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[3] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~2 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~2 .extended_lut = "off";
defparam \ShiftLeft0~2 .lut_mask = 64'h00E400E400E400E4;
defparam \ShiftLeft0~2 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[2] (
	.clk(clk_clk),
	.d(\ShiftLeft0~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[2]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[2] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[2] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[87]),
	.datac(!sink0_data[88]),
	.datad(!\in_size_reg[1]~q ),
	.datae(!\in_size_reg[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~3 .extended_lut = "off";
defparam \ShiftLeft0~3 .lut_mask = 64'hEA404040EA404040;
defparam \ShiftLeft0~3 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~4 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~4 .extended_lut = "off";
defparam \ShiftLeft0~4 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~4 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[1] (
	.clk(clk_clk),
	.d(\ShiftLeft0~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[1]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[1] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[1] .power_up = "low";

dffeas \int_byte_cnt_narrow_reg[0] (
	.clk(clk_clk),
	.d(\align_address_to_size|LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[0]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[0] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[0] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[0]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~3 (
	.dataa(!h2f_ARADDR_0),
	.datab(!sink0_data[69]),
	.datac(!sink0_data[68]),
	.datad(!out_data_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~3 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~3 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[0]~3 .shared_arith = "off";

dffeas \in_burstwrap_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[79]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[0]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[0] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[0] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[0]~0 (
	.dataa(!Selector13),
	.datab(!Selector6),
	.datac(!sink0_data[68]),
	.datad(!sink0_data[69]),
	.datae(!\new_burst_reg~q ),
	.dataf(!\d0_int_nxt_addr[0]~4_combout ),
	.datag(!\in_burstwrap_reg[0]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[0]~0 .extended_lut = "on";
defparam \nxt_addr[0]~0 .lut_mask = 64'h00000000F0F0FCA8;
defparam \nxt_addr[0]~0 .shared_arith = "off";

dffeas \int_nxt_addr_reg[0] (
	.clk(clk_clk),
	.d(\nxt_addr[0]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[0] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~4 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\Add0~13_sumout ),
	.datac(!\align_address_to_size|LessThan0~0_combout ),
	.datad(!\d0_int_nxt_addr[0]~3_combout ),
	.datae(!\int_nxt_addr_reg[0]~q ),
	.dataf(!\in_burstwrap_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~4 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~4 .lut_mask = 64'h0005AAAF2227AAAF;
defparam \d0_int_nxt_addr[0]~4 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[0] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[0]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[0] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[1]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[1]~q ),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \in_burstwrap_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[80]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[1]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[1] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[1] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[1]~4 (
	.dataa(!Selector12),
	.datab(!Selector5),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!\new_burst_reg~q ),
	.dataf(!\d0_int_nxt_addr[1]~2_combout ),
	.datag(!\in_burstwrap_reg[1]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[1]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[1]~4 .extended_lut = "on";
defparam \nxt_addr[1]~4 .lut_mask = 64'h00000000F0F0FAC8;
defparam \nxt_addr[1]~4 .shared_arith = "off";

dffeas \int_nxt_addr_reg[1] (
	.clk(clk_clk),
	.d(\nxt_addr[1]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[1] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~7 (
	.dataa(!h2f_ARADDR_1),
	.datab(!sink0_data[69]),
	.datac(!sink0_data[68]),
	.datad(!out_data_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~7 .extended_lut = "off";
defparam \d0_int_nxt_addr[1]~7 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[1]~7 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~2 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\Add0~9_sumout ),
	.datac(!\in_burstwrap_reg[1]~q ),
	.datad(!\int_nxt_addr_reg[1]~q ),
	.datae(!\ShiftLeft0~3_combout ),
	.dataf(!\d0_int_nxt_addr[1]~7_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~2 .extended_lut = "off";
defparam \d0_int_nxt_addr[1]~2 .lut_mask = 64'h02AA02AA02AA57FF;
defparam \d0_int_nxt_addr[1]~2 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[1] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[1]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[1] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_2),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[2]~q ),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[3]~q ),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

dffeas \in_burstwrap_reg[3] (
	.clk(clk_clk),
	.d(sink0_data[82]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[3]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[3] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[3] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[3]~12 (
	.dataa(!Selector10),
	.datab(!Selector3),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!\new_burst_reg~q ),
	.dataf(!\d0_int_nxt_addr[3]~0_combout ),
	.datag(!\in_burstwrap_reg[3]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[3]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[3]~12 .extended_lut = "on";
defparam \nxt_addr[3]~12 .lut_mask = 64'h00000000F0F0FAC8;
defparam \nxt_addr[3]~12 .shared_arith = "off";

dffeas \int_nxt_addr_reg[3] (
	.clk(clk_clk),
	.d(\nxt_addr[3]~12_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[3]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[3] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~5 (
	.dataa(!\Add0~1_sumout ),
	.datab(!\in_burstwrap_reg[3]~q ),
	.datac(!\int_nxt_addr_reg[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~5 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~5 .lut_mask = 64'hE0E0E0E0E0E0E0E0;
defparam \d0_int_nxt_addr[3]~5 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!h2f_ARADDR_3),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!base_address_3),
	.dataf(!\d0_int_nxt_addr[3]~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~0 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~0 .lut_mask = 64'hABABABFF01010155;
defparam \d0_int_nxt_addr[3]~0 .shared_arith = "off";

dffeas \in_burstwrap_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[81]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[2]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[2] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[2] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[2]~8 (
	.dataa(!Selector11),
	.datab(!Selector4),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!\new_burst_reg~q ),
	.dataf(!\d0_int_nxt_addr[2]~1_combout ),
	.datag(!\in_burstwrap_reg[2]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[2]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[2]~8 .extended_lut = "on";
defparam \nxt_addr[2]~8 .lut_mask = 64'h00000000F0F0FAC8;
defparam \nxt_addr[2]~8 .shared_arith = "off";

dffeas \int_nxt_addr_reg[2] (
	.clk(clk_clk),
	.d(\nxt_addr[2]~8_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[2]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~6 (
	.dataa(!\Add0~5_sumout ),
	.datab(!\in_burstwrap_reg[2]~q ),
	.datac(!\int_nxt_addr_reg[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~6 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~6 .lut_mask = 64'hE0E0E0E0E0E0E0E0;
defparam \d0_int_nxt_addr[2]~6 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!h2f_ARADDR_2),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!base_address_2),
	.dataf(!\d0_int_nxt_addr[2]~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~1 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~1 .lut_mask = 64'hABABABFF01010155;
defparam \d0_int_nxt_addr[2]~1 .shared_arith = "off";

dffeas in_eop_reg(
	.clk(clk_clk),
	.d(sink0_endofpacket),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_eop_reg~q ),
	.prn(vcc));
defparam in_eop_reg.is_wysiwyg = "true";
defparam in_eop_reg.power_up = "low";

endmodule

module spw_babasu_altera_merlin_address_alignment_11 (
	new_burst_reg,
	src_data_86,
	in_size_reg_0,
	ShiftLeft0,
	LessThan0)/* synthesis synthesis_greybox=0 */;
input 	new_burst_reg;
input 	src_data_86;
input 	in_size_reg_0;
input 	ShiftLeft0;
output 	LessThan0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!new_burst_reg),
	.datab(!src_data_86),
	.datac(!in_size_reg_0),
	.datad(!ShiftLeft0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan0),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h00E400E400E400E4;
defparam \LessThan0~0 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_burst_adapter_11 (
	h2f_ARADDR_0,
	h2f_ARADDR_1,
	h2f_ARADDR_2,
	h2f_ARADDR_3,
	h2f_ARBURST_0,
	h2f_ARBURST_1,
	h2f_ARID_0,
	h2f_ARID_1,
	h2f_ARID_2,
	h2f_ARID_3,
	h2f_ARID_4,
	h2f_ARID_5,
	h2f_ARID_6,
	h2f_ARID_7,
	h2f_ARID_8,
	h2f_ARID_9,
	h2f_ARID_10,
	h2f_ARID_11,
	h2f_ARLEN_0,
	Add5,
	Add51,
	in_ready_hold,
	saved_grant_1,
	stateST_COMP_TRANS,
	mem_used_1,
	in_data_reg_69,
	in_narrow_reg,
	cp_ready,
	cp_ready1,
	nxt_out_eop,
	out_valid_reg,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready,
	altera_reset_synchronizer_int_chain_out,
	Decoder1,
	Add2,
	Add21,
	Add22,
	Add23,
	nxt_in_ready1,
	src_valid,
	out_byte_cnt_reg_2,
	cp_ready2,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_6,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	Selector10,
	Selector101,
	Selector11,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	Selector12,
	src_payload,
	src_payload1,
	src_payload2,
	Selector13,
	nxt_out_burstwrap_1,
	nxt_addr_2,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARADDR_0;
input 	h2f_ARADDR_1;
input 	h2f_ARADDR_2;
input 	h2f_ARADDR_3;
input 	h2f_ARBURST_0;
input 	h2f_ARBURST_1;
input 	h2f_ARID_0;
input 	h2f_ARID_1;
input 	h2f_ARID_2;
input 	h2f_ARID_3;
input 	h2f_ARID_4;
input 	h2f_ARID_5;
input 	h2f_ARID_6;
input 	h2f_ARID_7;
input 	h2f_ARID_8;
input 	h2f_ARID_9;
input 	h2f_ARID_10;
input 	h2f_ARID_11;
input 	h2f_ARLEN_0;
input 	Add5;
input 	Add51;
input 	in_ready_hold;
input 	saved_grant_1;
output 	stateST_COMP_TRANS;
input 	mem_used_1;
output 	in_data_reg_69;
output 	in_narrow_reg;
input 	cp_ready;
input 	cp_ready1;
output 	nxt_out_eop;
output 	out_valid_reg;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready;
input 	altera_reset_synchronizer_int_chain_out;
input 	Decoder1;
input 	Add2;
input 	Add21;
input 	Add22;
input 	Add23;
output 	nxt_in_ready1;
input 	src_valid;
output 	out_byte_cnt_reg_2;
input 	cp_ready2;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_6;
output 	in_data_reg_105;
output 	in_data_reg_106;
output 	in_data_reg_107;
output 	in_data_reg_108;
output 	in_data_reg_109;
output 	in_data_reg_110;
output 	in_data_reg_111;
output 	in_data_reg_112;
output 	in_data_reg_113;
output 	in_data_reg_114;
output 	in_data_reg_115;
output 	in_data_reg_116;
input 	Selector10;
input 	Selector101;
input 	Selector11;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
input 	Selector12;
input 	src_payload;
input 	src_payload1;
input 	src_payload2;
input 	Selector13;
input 	nxt_out_burstwrap_1;
input 	nxt_addr_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



spw_babasu_altera_merlin_burst_adapter_13_1_11 \altera_merlin_burst_adapter_13_1.burst_adapter (
	.h2f_ARADDR_0(h2f_ARADDR_0),
	.h2f_ARADDR_1(h2f_ARADDR_1),
	.h2f_ARADDR_2(h2f_ARADDR_2),
	.h2f_ARADDR_3(h2f_ARADDR_3),
	.h2f_ARBURST_0(h2f_ARBURST_0),
	.h2f_ARBURST_1(h2f_ARBURST_1),
	.sink0_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,h2f_ARID_11,h2f_ARID_10,h2f_ARID_9,h2f_ARID_8,h2f_ARID_7,h2f_ARID_6,h2f_ARID_5,h2f_ARID_4,h2f_ARID_3,h2f_ARID_2,h2f_ARID_1,h2f_ARID_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_payload1,src_payload2,src_payload,gnd,gnd,gnd,
Selector101,Selector11,Selector12,Selector13,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,saved_grant_1,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.h2f_ARLEN_0(h2f_ARLEN_0),
	.Add5(Add5),
	.Add51(Add51),
	.in_ready_hold(in_ready_hold),
	.stateST_COMP_TRANS(stateST_COMP_TRANS),
	.mem_used_1(mem_used_1),
	.in_data_reg_69(in_data_reg_69),
	.in_narrow_reg1(in_narrow_reg),
	.cp_ready(cp_ready),
	.cp_ready1(cp_ready1),
	.nxt_out_eop(nxt_out_eop),
	.out_valid_reg1(out_valid_reg),
	.stateST_UNCOMP_WR_SUBBURST(stateST_UNCOMP_WR_SUBBURST),
	.nxt_in_ready(nxt_in_ready),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.Decoder1(Decoder1),
	.Add2(Add2),
	.Add21(Add21),
	.Add22(Add22),
	.Add23(Add23),
	.nxt_in_ready1(nxt_in_ready1),
	.src_valid(src_valid),
	.out_byte_cnt_reg_2(out_byte_cnt_reg_2),
	.cp_ready2(cp_ready2),
	.out_uncomp_byte_cnt_reg_3(out_uncomp_byte_cnt_reg_3),
	.out_uncomp_byte_cnt_reg_2(out_uncomp_byte_cnt_reg_2),
	.out_uncomp_byte_cnt_reg_4(out_uncomp_byte_cnt_reg_4),
	.out_uncomp_byte_cnt_reg_5(out_uncomp_byte_cnt_reg_5),
	.out_uncomp_byte_cnt_reg_6(out_uncomp_byte_cnt_reg_6),
	.in_data_reg_105(in_data_reg_105),
	.in_data_reg_106(in_data_reg_106),
	.in_data_reg_107(in_data_reg_107),
	.in_data_reg_108(in_data_reg_108),
	.in_data_reg_109(in_data_reg_109),
	.in_data_reg_110(in_data_reg_110),
	.in_data_reg_111(in_data_reg_111),
	.in_data_reg_112(in_data_reg_112),
	.in_data_reg_113(in_data_reg_113),
	.in_data_reg_114(in_data_reg_114),
	.in_data_reg_115(in_data_reg_115),
	.in_data_reg_116(in_data_reg_116),
	.Selector10(Selector10),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_3),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_2),
	.nxt_out_burstwrap_1(nxt_out_burstwrap_1),
	.nxt_addr_2(nxt_addr_2),
	.clk_clk(clk_clk));

endmodule

module spw_babasu_altera_merlin_burst_adapter_13_1_11 (
	h2f_ARADDR_0,
	h2f_ARADDR_1,
	h2f_ARADDR_2,
	h2f_ARADDR_3,
	h2f_ARBURST_0,
	h2f_ARBURST_1,
	sink0_data,
	h2f_ARLEN_0,
	Add5,
	Add51,
	in_ready_hold,
	stateST_COMP_TRANS,
	mem_used_1,
	in_data_reg_69,
	in_narrow_reg1,
	cp_ready,
	cp_ready1,
	nxt_out_eop,
	out_valid_reg1,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready,
	altera_reset_synchronizer_int_chain_out,
	Decoder1,
	Add2,
	Add21,
	Add22,
	Add23,
	nxt_in_ready1,
	src_valid,
	out_byte_cnt_reg_2,
	cp_ready2,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_6,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	Selector10,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	nxt_out_burstwrap_1,
	nxt_addr_2,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARADDR_0;
input 	h2f_ARADDR_1;
input 	h2f_ARADDR_2;
input 	h2f_ARADDR_3;
input 	h2f_ARBURST_0;
input 	h2f_ARBURST_1;
input 	[128:0] sink0_data;
input 	h2f_ARLEN_0;
input 	Add5;
input 	Add51;
input 	in_ready_hold;
output 	stateST_COMP_TRANS;
input 	mem_used_1;
output 	in_data_reg_69;
output 	in_narrow_reg1;
input 	cp_ready;
input 	cp_ready1;
output 	nxt_out_eop;
output 	out_valid_reg1;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready;
input 	altera_reset_synchronizer_int_chain_out;
input 	Decoder1;
input 	Add2;
input 	Add21;
input 	Add22;
input 	Add23;
output 	nxt_in_ready1;
input 	src_valid;
output 	out_byte_cnt_reg_2;
input 	cp_ready2;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_6;
output 	in_data_reg_105;
output 	in_data_reg_106;
output 	in_data_reg_107;
output 	in_data_reg_108;
output 	in_data_reg_109;
output 	in_data_reg_110;
output 	in_data_reg_111;
output 	in_data_reg_112;
output 	in_data_reg_113;
output 	in_data_reg_114;
output 	in_data_reg_115;
output 	in_data_reg_116;
input 	Selector10;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
input 	nxt_out_burstwrap_1;
input 	nxt_addr_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \align_address_to_size|LessThan0~0_combout ;
wire \align_address_to_size|LessThan0~1_combout ;
wire \nxt_uncomp_subburst_byte_cnt~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt[3]~1_combout ;
wire \nxt_uncomp_subburst_byte_cnt[4]~2_combout ;
wire \Add4~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt[5]~3_combout ;
wire \nxt_uncomp_subburst_byte_cnt[6]~4_combout ;
wire \nxt_uncomp_subburst_byte_cnt[2]~5_combout ;
wire \WideNor1~combout ;
wire \Selector2~1_combout ;
wire \load_next_out_cmd~combout ;
wire \state.ST_UNCOMP_TRANS~q ;
wire \Selector2~0_combout ;
wire \Selector0~0_combout ;
wire \state.ST_IDLE~q ;
wire \Selector1~0_combout ;
wire \Selector1~1_combout ;
wire \NON_PIPELINED_INPUTS.load_next_cmd~0_combout ;
wire \int_bytes_remaining_reg[3]~q ;
wire \d0_int_bytes_remaining[2]~4_combout ;
wire \int_bytes_remaining_reg[2]~q ;
wire \d0_int_bytes_remaining[3]~0_combout ;
wire \int_bytes_remaining_reg[4]~q ;
wire \Add1~0_combout ;
wire \d0_int_bytes_remaining[4]~1_combout ;
wire \int_bytes_remaining_reg[5]~q ;
wire \Add1~1_combout ;
wire \d0_int_bytes_remaining[5]~2_combout ;
wire \int_bytes_remaining_reg[6]~q ;
wire \d0_int_bytes_remaining[6]~3_combout ;
wire \new_burst_reg~0_combout ;
wire \new_burst_reg~q ;
wire \in_bytecount_reg_zero~0_combout ;
wire \in_bytecount_reg_zero~q ;
wire \nxt_out_valid~0_combout ;
wire \nxt_out_valid~1_combout ;
wire \Selector3~0_combout ;
wire \in_burstwrap_reg[3]~q ;
wire \nxt_addr[3]~0_combout ;
wire \nxt_addr[3]~combout ;
wire \int_nxt_addr_reg[3]~q ;
wire \in_size_reg[0]~q ;
wire \in_size_reg[2]~q ;
wire \in_size_reg[1]~q ;
wire \ShiftLeft0~0_combout ;
wire \ShiftLeft0~1_combout ;
wire \int_byte_cnt_narrow_reg[3]~q ;
wire \ShiftLeft0~2_combout ;
wire \int_byte_cnt_narrow_reg[2]~q ;
wire \in_burstwrap_reg[1]~q ;
wire \nxt_addr[1]~combout ;
wire \int_nxt_addr_reg[1]~q ;
wire \ShiftLeft0~3_combout ;
wire \int_byte_cnt_narrow_reg[1]~q ;
wire \int_byte_cnt_narrow_reg[0]~q ;
wire \Add0~13_sumout ;
wire \in_burstwrap_reg[0]~q ;
wire \nxt_addr[0]~combout ;
wire \int_nxt_addr_reg[0]~q ;
wire \d0_int_nxt_addr[0]~2_combout ;
wire \d0_int_nxt_addr[0]~3_combout ;
wire \int_nxt_addr_reg_dly[0]~q ;
wire \Add0~14 ;
wire \Add0~9_sumout ;
wire \d0_int_nxt_addr[1]~4_combout ;
wire \int_nxt_addr_reg_dly[1]~q ;
wire \Add0~10 ;
wire \Add0~6 ;
wire \Add0~1_sumout ;
wire \d0_int_nxt_addr[3]~0_combout ;
wire \in_burstwrap_reg[2]~q ;
wire \nxt_addr[2]~1_combout ;
wire \nxt_addr[2]~combout ;
wire \int_nxt_addr_reg[2]~q ;
wire \Add0~5_sumout ;
wire \d0_int_nxt_addr[2]~1_combout ;


spw_babasu_altera_merlin_address_alignment_12 align_address_to_size(
	.new_burst_reg(\new_burst_reg~q ),
	.src_payload(sink0_data[86]),
	.in_size_reg_0(\in_size_reg[0]~q ),
	.src_payload1(sink0_data[88]),
	.in_size_reg_2(\in_size_reg[2]~q ),
	.src_payload2(sink0_data[87]),
	.in_size_reg_1(\in_size_reg[1]~q ),
	.LessThan0(\align_address_to_size|LessThan0~0_combout ),
	.LessThan01(\align_address_to_size|LessThan0~1_combout ));

dffeas \state.ST_COMP_TRANS (
	.clk(clk_clk),
	.d(\Selector1~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_COMP_TRANS),
	.prn(vcc));
defparam \state.ST_COMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_COMP_TRANS .power_up = "low";

dffeas \in_data_reg[69] (
	.clk(clk_clk),
	.d(sink0_data[69]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_69),
	.prn(vcc));
defparam \in_data_reg[69] .is_wysiwyg = "true";
defparam \in_data_reg[69] .power_up = "low";

dffeas in_narrow_reg(
	.clk(clk_clk),
	.d(Decoder1),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_narrow_reg1),
	.prn(vcc));
defparam in_narrow_reg.is_wysiwyg = "true";
defparam in_narrow_reg.power_up = "low";

cyclonev_lcell_comb \nxt_out_eop~0 (
	.dataa(!in_data_reg_69),
	.datab(!stateST_COMP_TRANS),
	.datac(!\new_burst_reg~q ),
	.datad(!mem_used_1),
	.datae(!cp_ready),
	.dataf(!\in_bytecount_reg_zero~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_out_eop),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_eop~0 .extended_lut = "off";
defparam \nxt_out_eop~0 .lut_mask = 64'h4444474477774777;
defparam \nxt_out_eop~0 .shared_arith = "off";

dffeas out_valid_reg(
	.clk(clk_clk),
	.d(\nxt_out_valid~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_valid_reg1),
	.prn(vcc));
defparam out_valid_reg.is_wysiwyg = "true";
defparam out_valid_reg.power_up = "low";

dffeas \state.ST_UNCOMP_WR_SUBBURST (
	.clk(clk_clk),
	.d(\Selector3~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_UNCOMP_WR_SUBBURST),
	.prn(vcc));
defparam \state.ST_UNCOMP_WR_SUBBURST .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_WR_SUBBURST .power_up = "low";

cyclonev_lcell_comb \nxt_in_ready~0 (
	.dataa(!in_ready_hold),
	.datab(!stateST_COMP_TRANS),
	.datac(!mem_used_1),
	.datad(!cp_ready),
	.datae(!out_valid_reg1),
	.dataf(!\Selector2~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~0 .extended_lut = "off";
defparam \nxt_in_ready~0 .lut_mask = 64'h0000FF3F8888BBBB;
defparam \nxt_in_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_in_ready~1 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!cp_ready1),
	.datac(!nxt_out_eop),
	.datad(!nxt_in_ready),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~1 .extended_lut = "off";
defparam \nxt_in_ready~1 .lut_mask = 64'h00FE00FE00FE00FE;
defparam \nxt_in_ready~1 .shared_arith = "off";

dffeas \out_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[3] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[3]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_3),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[3] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[3] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[2]~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[4] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[4]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_4),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[4] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[4] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[5] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[5]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_5),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[5] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[5] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[6] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[6]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_6),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[6] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[6] .power_up = "low";

dffeas \in_data_reg[105] (
	.clk(clk_clk),
	.d(sink0_data[105]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_105),
	.prn(vcc));
defparam \in_data_reg[105] .is_wysiwyg = "true";
defparam \in_data_reg[105] .power_up = "low";

dffeas \in_data_reg[106] (
	.clk(clk_clk),
	.d(sink0_data[106]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_106),
	.prn(vcc));
defparam \in_data_reg[106] .is_wysiwyg = "true";
defparam \in_data_reg[106] .power_up = "low";

dffeas \in_data_reg[107] (
	.clk(clk_clk),
	.d(sink0_data[107]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_107),
	.prn(vcc));
defparam \in_data_reg[107] .is_wysiwyg = "true";
defparam \in_data_reg[107] .power_up = "low";

dffeas \in_data_reg[108] (
	.clk(clk_clk),
	.d(sink0_data[108]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_108),
	.prn(vcc));
defparam \in_data_reg[108] .is_wysiwyg = "true";
defparam \in_data_reg[108] .power_up = "low";

dffeas \in_data_reg[109] (
	.clk(clk_clk),
	.d(sink0_data[109]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_109),
	.prn(vcc));
defparam \in_data_reg[109] .is_wysiwyg = "true";
defparam \in_data_reg[109] .power_up = "low";

dffeas \in_data_reg[110] (
	.clk(clk_clk),
	.d(sink0_data[110]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_110),
	.prn(vcc));
defparam \in_data_reg[110] .is_wysiwyg = "true";
defparam \in_data_reg[110] .power_up = "low";

dffeas \in_data_reg[111] (
	.clk(clk_clk),
	.d(sink0_data[111]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_111),
	.prn(vcc));
defparam \in_data_reg[111] .is_wysiwyg = "true";
defparam \in_data_reg[111] .power_up = "low";

dffeas \in_data_reg[112] (
	.clk(clk_clk),
	.d(sink0_data[112]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_112),
	.prn(vcc));
defparam \in_data_reg[112] .is_wysiwyg = "true";
defparam \in_data_reg[112] .power_up = "low";

dffeas \in_data_reg[113] (
	.clk(clk_clk),
	.d(sink0_data[113]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_113),
	.prn(vcc));
defparam \in_data_reg[113] .is_wysiwyg = "true";
defparam \in_data_reg[113] .power_up = "low";

dffeas \in_data_reg[114] (
	.clk(clk_clk),
	.d(sink0_data[114]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_114),
	.prn(vcc));
defparam \in_data_reg[114] .is_wysiwyg = "true";
defparam \in_data_reg[114] .power_up = "low";

dffeas \in_data_reg[115] (
	.clk(clk_clk),
	.d(sink0_data[115]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_115),
	.prn(vcc));
defparam \in_data_reg[115] .is_wysiwyg = "true";
defparam \in_data_reg[115] .power_up = "low";

dffeas \in_data_reg[116] (
	.clk(clk_clk),
	.d(sink0_data[116]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_116),
	.prn(vcc));
defparam \in_data_reg[116] .is_wysiwyg = "true";
defparam \in_data_reg[116] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[3] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[3]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_3),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[3] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[2] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[2]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_2),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[2] .power_up = "low";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt~0 (
	.dataa(!cp_ready1),
	.datab(!out_valid_reg1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt~0 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt~0 .lut_mask = 64'h1111111111111111;
defparam \nxt_uncomp_subburst_byte_cnt~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[3]~1 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!out_uncomp_byte_cnt_reg_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[3]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[3]~1 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[3]~1 .lut_mask = 64'h0FE40F4E0FE40F4E;
defparam \nxt_uncomp_subburst_byte_cnt[3]~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[4]~2 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!out_uncomp_byte_cnt_reg_2),
	.dataf(!out_uncomp_byte_cnt_reg_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[4]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[4]~2 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[4]~2 .lut_mask = 64'h00E40044FF4EFFEE;
defparam \nxt_uncomp_subburst_byte_cnt[4]~2 .shared_arith = "off";

cyclonev_lcell_comb \Add4~0 (
	.dataa(!out_uncomp_byte_cnt_reg_3),
	.datab(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datac(!out_uncomp_byte_cnt_reg_2),
	.datad(!out_uncomp_byte_cnt_reg_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add4~0 .extended_lut = "off";
defparam \Add4~0 .lut_mask = 64'h2000200020002000;
defparam \Add4~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[5]~3 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_5),
	.datae(!\Add4~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[5]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[5]~3 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[5]~3 .lut_mask = 64'h04FEAE5404FEAE54;
defparam \nxt_uncomp_subburst_byte_cnt[5]~3 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[6]~4 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_5),
	.datae(!\Add4~0_combout ),
	.dataf(!out_uncomp_byte_cnt_reg_6),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[6]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[6]~4 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[6]~4 .lut_mask = 64'h0404AE04FEFE54FE;
defparam \nxt_uncomp_subburst_byte_cnt[6]~4 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[2]~5 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[2]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[2]~5 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[2]~5 .lut_mask = 64'h0EF40EF40EF40EF4;
defparam \nxt_uncomp_subburst_byte_cnt[2]~5 .shared_arith = "off";

cyclonev_lcell_comb WideNor1(
	.dataa(!\nxt_uncomp_subburst_byte_cnt[3]~1_combout ),
	.datab(!\nxt_uncomp_subburst_byte_cnt[4]~2_combout ),
	.datac(!\nxt_uncomp_subburst_byte_cnt[5]~3_combout ),
	.datad(!\nxt_uncomp_subburst_byte_cnt[6]~4_combout ),
	.datae(!\nxt_uncomp_subburst_byte_cnt[2]~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideNor1.extended_lut = "off";
defparam WideNor1.lut_mask = 64'h8000000080000000;
defparam WideNor1.shared_arith = "off";

cyclonev_lcell_comb \Selector2~1 (
	.dataa(!nxt_out_eop),
	.datab(!\Selector2~0_combout ),
	.datac(!\WideNor1~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~1 .extended_lut = "off";
defparam \Selector2~1 .lut_mask = 64'h0808080808080808;
defparam \Selector2~1 .shared_arith = "off";

cyclonev_lcell_comb load_next_out_cmd(
	.dataa(!mem_used_1),
	.datab(!cp_ready),
	.datac(!out_valid_reg1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\load_next_out_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam load_next_out_cmd.extended_lut = "off";
defparam load_next_out_cmd.lut_mask = 64'hF2F2F2F2F2F2F2F2;
defparam load_next_out_cmd.shared_arith = "off";

dffeas \state.ST_UNCOMP_TRANS (
	.clk(clk_clk),
	.d(\Selector2~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_UNCOMP_TRANS~q ),
	.prn(vcc));
defparam \state.ST_UNCOMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_TRANS .power_up = "low";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'h8888888888888888;
defparam \Selector2~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!in_ready_hold),
	.datab(!nxt_out_eop),
	.datac(!src_valid),
	.datad(!\state.ST_IDLE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'h05CD05CD05CD05CD;
defparam \Selector0~0 .shared_arith = "off";

dffeas \state.ST_IDLE (
	.clk(clk_clk),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_IDLE~q ),
	.prn(vcc));
defparam \state.ST_IDLE .is_wysiwyg = "true";
defparam \state.ST_IDLE .power_up = "low";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!sink0_data[69]),
	.datab(!nxt_out_eop),
	.datac(!\Selector2~0_combout ),
	.datad(!\state.ST_IDLE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'h5510551055105510;
defparam \Selector1~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~1 (
	.dataa(!in_ready_hold),
	.datab(!stateST_COMP_TRANS),
	.datac(!nxt_out_eop),
	.datad(!src_valid),
	.datae(!\Selector1~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~1 .extended_lut = "off";
defparam \Selector1~1 .lut_mask = 64'h3031307530313075;
defparam \Selector1~1 .shared_arith = "off";

cyclonev_lcell_comb \NON_PIPELINED_INPUTS.load_next_cmd~0 (
	.dataa(!in_ready_hold),
	.datab(!nxt_in_ready1),
	.datac(!src_valid),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \NON_PIPELINED_INPUTS.load_next_cmd~0 .extended_lut = "off";
defparam \NON_PIPELINED_INPUTS.load_next_cmd~0 .lut_mask = 64'h0404040404040404;
defparam \NON_PIPELINED_INPUTS.load_next_cmd~0 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[3] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[3]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[3]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[3] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[3] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[2]~4 (
	.dataa(!h2f_ARLEN_0),
	.datab(!sink0_data[69]),
	.datac(!\new_burst_reg~q ),
	.datad(!out_byte_cnt_reg_2),
	.datae(!\int_bytes_remaining_reg[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[2]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[2]~4 .extended_lut = "off";
defparam \d0_int_bytes_remaining[2]~4 .lut_mask = 64'h02F2F20202F2F202;
defparam \d0_int_bytes_remaining[2]~4 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[2] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[2]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[2]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[2] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[3]~0 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!Add2),
	.datad(!\int_bytes_remaining_reg[3]~q ),
	.datae(!out_byte_cnt_reg_2),
	.dataf(!\int_bytes_remaining_reg[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[3]~0 .extended_lut = "off";
defparam \d0_int_bytes_remaining[3]~0 .lut_mask = 64'h01CDCD0101CD01CD;
defparam \d0_int_bytes_remaining[3]~0 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[4] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[4]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[4]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[4] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[4] .power_up = "low";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!\int_bytes_remaining_reg[3]~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\int_bytes_remaining_reg[2]~q ),
	.datad(!\int_bytes_remaining_reg[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'hDF20DF20DF20DF20;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[4]~1 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!Add21),
	.datad(!\Add1~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[4]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[4]~1 .extended_lut = "off";
defparam \d0_int_bytes_remaining[4]~1 .lut_mask = 64'hCD01CD01CD01CD01;
defparam \d0_int_bytes_remaining[4]~1 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[5] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[5]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[5]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[5] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[5] .power_up = "low";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!\int_bytes_remaining_reg[3]~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\int_bytes_remaining_reg[2]~q ),
	.datad(!\int_bytes_remaining_reg[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h2000200020002000;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[5]~2 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!Add22),
	.datad(!\int_bytes_remaining_reg[5]~q ),
	.datae(!\Add1~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[5]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[5]~2 .extended_lut = "off";
defparam \d0_int_bytes_remaining[5]~2 .lut_mask = 64'h01CDCD0101CDCD01;
defparam \d0_int_bytes_remaining[5]~2 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[6] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[6]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[6]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[6] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[6] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[6]~3 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!Add23),
	.datad(!\int_bytes_remaining_reg[5]~q ),
	.datae(!\Add1~1_combout ),
	.dataf(!\int_bytes_remaining_reg[6]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[6]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[6]~3 .extended_lut = "off";
defparam \d0_int_bytes_remaining[6]~3 .lut_mask = 64'h0101CD01CDCD01CD;
defparam \d0_int_bytes_remaining[6]~3 .shared_arith = "off";

cyclonev_lcell_comb \new_burst_reg~0 (
	.dataa(!\Selector1~1_combout ),
	.datab(!\d0_int_bytes_remaining[3]~0_combout ),
	.datac(!\d0_int_bytes_remaining[4]~1_combout ),
	.datad(!\d0_int_bytes_remaining[5]~2_combout ),
	.datae(!\d0_int_bytes_remaining[6]~3_combout ),
	.dataf(!\d0_int_bytes_remaining[2]~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\new_burst_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \new_burst_reg~0 .extended_lut = "off";
defparam \new_burst_reg~0 .lut_mask = 64'hAAAAAAAAEAAAAAAA;
defparam \new_burst_reg~0 .shared_arith = "off";

dffeas new_burst_reg(
	.clk(clk_clk),
	.d(\new_burst_reg~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\new_burst_reg~q ),
	.prn(vcc));
defparam new_burst_reg.is_wysiwyg = "true";
defparam new_burst_reg.power_up = "low";

cyclonev_lcell_comb \in_bytecount_reg_zero~0 (
	.dataa(!sink0_data[69]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\in_bytecount_reg_zero~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \in_bytecount_reg_zero~0 .extended_lut = "off";
defparam \in_bytecount_reg_zero~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \in_bytecount_reg_zero~0 .shared_arith = "off";

dffeas in_bytecount_reg_zero(
	.clk(clk_clk),
	.d(\in_bytecount_reg_zero~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_bytecount_reg_zero~q ),
	.prn(vcc));
defparam in_bytecount_reg_zero.is_wysiwyg = "true";
defparam in_bytecount_reg_zero.power_up = "low";

cyclonev_lcell_comb \nxt_out_valid~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!mem_used_1),
	.datac(!\in_bytecount_reg_zero~q ),
	.datad(!cp_ready2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_valid~0 .extended_lut = "off";
defparam \nxt_out_valid~0 .lut_mask = 64'hF0B8F0B8F0B8F0B8;
defparam \nxt_out_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_out_valid~1 (
	.dataa(!in_ready_hold),
	.datab(!stateST_COMP_TRANS),
	.datac(!src_valid),
	.datad(!\nxt_out_valid~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_valid~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_valid~1 .extended_lut = "off";
defparam \nxt_out_valid~1 .lut_mask = 64'h0537053705370537;
defparam \nxt_out_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~0 (
	.dataa(!nxt_out_eop),
	.datab(!\Selector2~0_combout ),
	.datac(!\WideNor1~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'h8080808080808080;
defparam \Selector3~0 .shared_arith = "off";

dffeas \in_burstwrap_reg[3] (
	.clk(clk_clk),
	.d(sink0_data[82]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_burstwrap_reg[3]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[3] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[3] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[3]~0 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!\in_burstwrap_reg[3]~q ),
	.datad(!\d0_int_nxt_addr[3]~0_combout ),
	.datae(!h2f_ARBURST_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[3]~0 .extended_lut = "off";
defparam \nxt_addr[3]~0 .lut_mask = 64'h00F300E200F300E2;
defparam \nxt_addr[3]~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_addr[3] (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!h2f_ARBURST_1),
	.datad(!Add5),
	.datae(!Selector10),
	.dataf(!\nxt_addr[3]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[3] .extended_lut = "off";
defparam \nxt_addr[3] .lut_mask = 64'h00000000FEEEFFEF;
defparam \nxt_addr[3] .shared_arith = "off";

dffeas \int_nxt_addr_reg[3] (
	.clk(clk_clk),
	.d(\nxt_addr[3]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[3]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[3] .power_up = "low";

dffeas \in_size_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[86]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_size_reg[0]~q ),
	.prn(vcc));
defparam \in_size_reg[0] .is_wysiwyg = "true";
defparam \in_size_reg[0] .power_up = "low";

dffeas \in_size_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[88]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_size_reg[2]~q ),
	.prn(vcc));
defparam \in_size_reg[2] .is_wysiwyg = "true";
defparam \in_size_reg[2] .power_up = "low";

dffeas \in_size_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[87]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_size_reg[1]~q ),
	.prn(vcc));
defparam \in_size_reg[1] .is_wysiwyg = "true";
defparam \in_size_reg[1] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[88]),
	.datac(!\in_size_reg[2]~q ),
	.datad(!sink0_data[87]),
	.datae(!\in_size_reg[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~0 .extended_lut = "off";
defparam \ShiftLeft0~0 .lut_mask = 64'h0044A0E40044A0E4;
defparam \ShiftLeft0~0 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~1 .extended_lut = "off";
defparam \ShiftLeft0~1 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~1 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[3] (
	.clk(clk_clk),
	.d(\ShiftLeft0~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[3]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[3] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[3] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~2 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~2 .extended_lut = "off";
defparam \ShiftLeft0~2 .lut_mask = 64'h00E400E400E400E4;
defparam \ShiftLeft0~2 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[2] (
	.clk(clk_clk),
	.d(\ShiftLeft0~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[2]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[2] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[2] .power_up = "low";

dffeas \in_burstwrap_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[80]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_burstwrap_reg[1]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[1] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[1] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[1] (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!\in_burstwrap_reg[1]~q ),
	.datad(!\d0_int_nxt_addr[1]~4_combout ),
	.datae(!nxt_out_burstwrap_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[1] .extended_lut = "off";
defparam \nxt_addr[1] .lut_mask = 64'h00E200F300E200F3;
defparam \nxt_addr[1] .shared_arith = "off";

dffeas \int_nxt_addr_reg[1] (
	.clk(clk_clk),
	.d(\nxt_addr[1]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[1] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\align_address_to_size|LessThan0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~3 .extended_lut = "off";
defparam \ShiftLeft0~3 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~3 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[1] (
	.clk(clk_clk),
	.d(\ShiftLeft0~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[1]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[1] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[1] .power_up = "low";

dffeas \int_byte_cnt_narrow_reg[0] (
	.clk(clk_clk),
	.d(\align_address_to_size|LessThan0~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[0]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[0] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[0] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[0]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \in_burstwrap_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[79]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_burstwrap_reg[0]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[0] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[0] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[0] (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!sink0_data[79]),
	.datad(!\in_burstwrap_reg[0]~q ),
	.datae(!\d0_int_nxt_addr[0]~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[0] .extended_lut = "off";
defparam \nxt_addr[0] .lut_mask = 64'h0000FE320000FE32;
defparam \nxt_addr[0] .shared_arith = "off";

dffeas \int_nxt_addr_reg[0] (
	.clk(clk_clk),
	.d(\nxt_addr[0]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[0] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~2 (
	.dataa(!\Add0~13_sumout ),
	.datab(!\int_nxt_addr_reg[0]~q ),
	.datac(!\in_burstwrap_reg[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~2 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~2 .lut_mask = 64'hC8C8C8C8C8C8C8C8;
defparam \d0_int_nxt_addr[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~3 (
	.dataa(!h2f_ARADDR_0),
	.datab(!sink0_data[69]),
	.datac(!\new_burst_reg~q ),
	.datad(!\align_address_to_size|LessThan0~1_combout ),
	.datae(!\d0_int_nxt_addr[0]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~3 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~3 .lut_mask = 64'hF0F10001F0F10001;
defparam \d0_int_nxt_addr[0]~3 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[0] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[0]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[0] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[1]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[1]~q ),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~4 (
	.dataa(!\int_nxt_addr_reg[1]~q ),
	.datab(!\Add0~9_sumout ),
	.datac(!sink0_data[69]),
	.datad(!Decoder1),
	.datae(!\new_burst_reg~q ),
	.dataf(!h2f_ARADDR_1),
	.datag(!\in_burstwrap_reg[1]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~4 .extended_lut = "on";
defparam \d0_int_nxt_addr[1]~4 .lut_mask = 64'h575700005757000F;
defparam \d0_int_nxt_addr[1]~4 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[1] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[1]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[1] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_2),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[2]~q ),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[3]~q ),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~0 (
	.dataa(!h2f_ARADDR_3),
	.datab(!sink0_data[69]),
	.datac(!\new_burst_reg~q ),
	.datad(!\int_nxt_addr_reg[3]~q ),
	.datae(!\in_burstwrap_reg[3]~q ),
	.dataf(!\Add0~1_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~0 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~0 .lut_mask = 64'h01F101F101F1F1F1;
defparam \d0_int_nxt_addr[3]~0 .shared_arith = "off";

dffeas \in_burstwrap_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[81]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_burstwrap_reg[2]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[2] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[2] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[2]~1 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!\in_burstwrap_reg[2]~q ),
	.datad(!\d0_int_nxt_addr[2]~1_combout ),
	.datae(!h2f_ARBURST_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[2]~1 .extended_lut = "off";
defparam \nxt_addr[2]~1 .lut_mask = 64'h00F300E200F300E2;
defparam \nxt_addr[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_addr[2] (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!h2f_ARBURST_1),
	.datad(!Add51),
	.datae(!\nxt_addr[2]~1_combout ),
	.dataf(!nxt_addr_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[2] .extended_lut = "off";
defparam \nxt_addr[2] .lut_mask = 64'h0000FEEE0000FFEF;
defparam \nxt_addr[2] .shared_arith = "off";

dffeas \int_nxt_addr_reg[2] (
	.clk(clk_clk),
	.d(\nxt_addr[2]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[2]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~1 (
	.dataa(!h2f_ARADDR_2),
	.datab(!sink0_data[69]),
	.datac(!\new_burst_reg~q ),
	.datad(!\int_nxt_addr_reg[2]~q ),
	.datae(!\in_burstwrap_reg[2]~q ),
	.dataf(!\Add0~5_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~1 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~1 .lut_mask = 64'h01F101F101F1F1F1;
defparam \d0_int_nxt_addr[2]~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_address_alignment_12 (
	new_burst_reg,
	src_payload,
	in_size_reg_0,
	src_payload1,
	in_size_reg_2,
	src_payload2,
	in_size_reg_1,
	LessThan0,
	LessThan01)/* synthesis synthesis_greybox=0 */;
input 	new_burst_reg;
input 	src_payload;
input 	in_size_reg_0;
input 	src_payload1;
input 	in_size_reg_2;
input 	src_payload2;
input 	in_size_reg_1;
output 	LessThan0;
output 	LessThan01;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!new_burst_reg),
	.datab(!src_payload1),
	.datac(!in_size_reg_2),
	.datad(!src_payload2),
	.datae(!in_size_reg_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan0),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'hE4A04400E4A04400;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~1 (
	.dataa(!new_burst_reg),
	.datab(!src_payload),
	.datac(!in_size_reg_0),
	.datad(!LessThan0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan01),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~1 .extended_lut = "off";
defparam \LessThan0~1 .lut_mask = 64'h00E400E400E400E4;
defparam \LessThan0~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_burst_adapter_12 (
	h2f_ARADDR_0,
	h2f_ARADDR_1,
	h2f_ARADDR_2,
	h2f_ARADDR_3,
	h2f_ARLEN_0,
	nxt_in_ready,
	in_ready_hold,
	stateST_COMP_TRANS,
	out_valid_reg,
	in_narrow_reg,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	in_data_reg_68,
	cp_ready,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready1,
	saved_grant_1,
	Equal13,
	saved_grant_0,
	altera_reset_synchronizer_int_chain_out,
	in_data_reg_0,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	in_data_reg_1,
	in_data_reg_2,
	in_data_reg_3,
	in_data_reg_4,
	in_data_reg_5,
	in_data_reg_6,
	in_data_reg_7,
	Add2,
	Add21,
	Add22,
	Add23,
	write_cp_data_77,
	write_cp_data_78,
	write_cp_data_75,
	write_cp_data_74,
	write_cp_data_76,
	WideNor0,
	nxt_out_eop,
	Equal14,
	src14_valid,
	src_valid,
	cp_ready1,
	in_data_reg_69,
	src_data_87,
	src_data_88,
	src_valid1,
	src_data_35,
	src_data_34,
	src_data_33,
	src_data_32,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_6,
	src_payload_0,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	Selector3,
	Selector10,
	base_address_3,
	Selector4,
	Selector11,
	base_address_2,
	src_payload,
	src_data_82,
	src_data_81,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_data_105,
	src_data_106,
	src_data_107,
	src_data_108,
	src_data_109,
	src_data_110,
	src_data_111,
	src_data_112,
	src_data_113,
	src_data_114,
	src_data_115,
	src_data_116,
	src_data_86,
	Selector5,
	Selector12,
	out_data_1,
	src_data_80,
	out_data_0,
	Selector6,
	Selector13,
	src_data_79,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARADDR_0;
input 	h2f_ARADDR_1;
input 	h2f_ARADDR_2;
input 	h2f_ARADDR_3;
input 	h2f_ARLEN_0;
output 	nxt_in_ready;
input 	in_ready_hold;
output 	stateST_COMP_TRANS;
output 	out_valid_reg;
output 	in_narrow_reg;
output 	in_byteen_reg_3;
output 	in_byteen_reg_2;
output 	in_byteen_reg_1;
output 	in_byteen_reg_0;
output 	in_data_reg_68;
input 	cp_ready;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready1;
input 	saved_grant_1;
input 	Equal13;
input 	saved_grant_0;
input 	altera_reset_synchronizer_int_chain_out;
output 	in_data_reg_0;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
output 	in_data_reg_1;
output 	in_data_reg_2;
output 	in_data_reg_3;
output 	in_data_reg_4;
output 	in_data_reg_5;
output 	in_data_reg_6;
output 	in_data_reg_7;
input 	Add2;
input 	Add21;
input 	Add22;
input 	Add23;
input 	write_cp_data_77;
input 	write_cp_data_78;
input 	write_cp_data_75;
input 	write_cp_data_74;
input 	write_cp_data_76;
input 	WideNor0;
output 	nxt_out_eop;
input 	Equal14;
input 	src14_valid;
input 	src_valid;
input 	cp_ready1;
output 	in_data_reg_69;
input 	src_data_87;
input 	src_data_88;
input 	src_valid1;
input 	src_data_35;
input 	src_data_34;
input 	src_data_33;
input 	src_data_32;
output 	out_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_6;
input 	src_payload_0;
output 	in_data_reg_105;
output 	in_data_reg_106;
output 	in_data_reg_107;
output 	in_data_reg_108;
output 	in_data_reg_109;
output 	in_data_reg_110;
output 	in_data_reg_111;
output 	in_data_reg_112;
output 	in_data_reg_113;
output 	in_data_reg_114;
output 	in_data_reg_115;
output 	in_data_reg_116;
input 	Selector3;
input 	Selector10;
input 	base_address_3;
input 	Selector4;
input 	Selector11;
input 	base_address_2;
input 	src_payload;
input 	src_data_82;
input 	src_data_81;
input 	src_payload1;
input 	src_payload2;
input 	src_payload3;
input 	src_payload4;
input 	src_payload5;
input 	src_payload6;
input 	src_payload7;
input 	src_data_105;
input 	src_data_106;
input 	src_data_107;
input 	src_data_108;
input 	src_data_109;
input 	src_data_110;
input 	src_data_111;
input 	src_data_112;
input 	src_data_113;
input 	src_data_114;
input 	src_data_115;
input 	src_data_116;
input 	src_data_86;
input 	Selector5;
input 	Selector12;
input 	out_data_1;
input 	src_data_80;
input 	out_data_0;
input 	Selector6;
input 	Selector13;
input 	src_data_79;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



spw_babasu_altera_merlin_burst_adapter_13_1_12 \altera_merlin_burst_adapter_13_1.burst_adapter (
	.h2f_ARADDR_0(h2f_ARADDR_0),
	.h2f_ARADDR_1(h2f_ARADDR_1),
	.h2f_ARADDR_2(h2f_ARADDR_2),
	.h2f_ARADDR_3(h2f_ARADDR_3),
	.h2f_ARLEN_0(h2f_ARLEN_0),
	.nxt_in_ready(nxt_in_ready),
	.in_ready_hold(in_ready_hold),
	.stateST_COMP_TRANS(stateST_COMP_TRANS),
	.out_valid_reg1(out_valid_reg),
	.in_narrow_reg1(in_narrow_reg),
	.in_byteen_reg_3(in_byteen_reg_3),
	.in_byteen_reg_2(in_byteen_reg_2),
	.in_byteen_reg_1(in_byteen_reg_1),
	.in_byteen_reg_0(in_byteen_reg_0),
	.in_data_reg_68(in_data_reg_68),
	.cp_ready(cp_ready),
	.stateST_UNCOMP_WR_SUBBURST(stateST_UNCOMP_WR_SUBBURST),
	.nxt_in_ready1(nxt_in_ready1),
	.sink0_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_116,src_data_115,src_data_114,src_data_113,src_data_112,src_data_111,src_data_110,src_data_109,src_data_108,src_data_107,src_data_106,src_data_105,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_88,src_data_87,
src_data_86,gnd,gnd,gnd,src_data_82,src_data_81,src_data_80,src_data_79,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,saved_grant_1,saved_grant_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_35,src_data_34,src_data_33,
src_data_32,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_payload7,src_payload6,src_payload5,src_payload4,src_payload3,src_payload2,src_payload1,src_payload}),
	.Equal13(Equal13),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.in_data_reg_0(in_data_reg_0),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_3),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_2),
	.in_data_reg_1(in_data_reg_1),
	.in_data_reg_2(in_data_reg_2),
	.in_data_reg_3(in_data_reg_3),
	.in_data_reg_4(in_data_reg_4),
	.in_data_reg_5(in_data_reg_5),
	.in_data_reg_6(in_data_reg_6),
	.in_data_reg_7(in_data_reg_7),
	.Add2(Add2),
	.Add21(Add21),
	.Add22(Add22),
	.Add23(Add23),
	.write_cp_data_77(write_cp_data_77),
	.write_cp_data_78(write_cp_data_78),
	.write_cp_data_75(write_cp_data_75),
	.write_cp_data_74(write_cp_data_74),
	.write_cp_data_76(write_cp_data_76),
	.WideNor0(WideNor0),
	.nxt_out_eop(nxt_out_eop),
	.Equal14(Equal14),
	.src14_valid(src14_valid),
	.src_valid(src_valid),
	.cp_ready1(cp_ready1),
	.in_data_reg_69(in_data_reg_69),
	.src_valid1(src_valid1),
	.out_byte_cnt_reg_2(out_byte_cnt_reg_2),
	.out_uncomp_byte_cnt_reg_5(out_uncomp_byte_cnt_reg_5),
	.out_uncomp_byte_cnt_reg_4(out_uncomp_byte_cnt_reg_4),
	.out_uncomp_byte_cnt_reg_3(out_uncomp_byte_cnt_reg_3),
	.out_uncomp_byte_cnt_reg_2(out_uncomp_byte_cnt_reg_2),
	.out_uncomp_byte_cnt_reg_6(out_uncomp_byte_cnt_reg_6),
	.sink0_endofpacket(src_payload_0),
	.in_data_reg_105(in_data_reg_105),
	.in_data_reg_106(in_data_reg_106),
	.in_data_reg_107(in_data_reg_107),
	.in_data_reg_108(in_data_reg_108),
	.in_data_reg_109(in_data_reg_109),
	.in_data_reg_110(in_data_reg_110),
	.in_data_reg_111(in_data_reg_111),
	.in_data_reg_112(in_data_reg_112),
	.in_data_reg_113(in_data_reg_113),
	.in_data_reg_114(in_data_reg_114),
	.in_data_reg_115(in_data_reg_115),
	.in_data_reg_116(in_data_reg_116),
	.Selector3(Selector3),
	.Selector10(Selector10),
	.base_address_3(base_address_3),
	.Selector4(Selector4),
	.Selector11(Selector11),
	.base_address_2(base_address_2),
	.Selector5(Selector5),
	.Selector12(Selector12),
	.out_data_1(out_data_1),
	.out_data_0(out_data_0),
	.Selector6(Selector6),
	.Selector13(Selector13),
	.clk_clk(clk_clk));

endmodule

module spw_babasu_altera_merlin_burst_adapter_13_1_12 (
	h2f_ARADDR_0,
	h2f_ARADDR_1,
	h2f_ARADDR_2,
	h2f_ARADDR_3,
	h2f_ARLEN_0,
	nxt_in_ready,
	in_ready_hold,
	stateST_COMP_TRANS,
	out_valid_reg1,
	in_narrow_reg1,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	in_data_reg_68,
	cp_ready,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready1,
	sink0_data,
	Equal13,
	altera_reset_synchronizer_int_chain_out,
	in_data_reg_0,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	in_data_reg_1,
	in_data_reg_2,
	in_data_reg_3,
	in_data_reg_4,
	in_data_reg_5,
	in_data_reg_6,
	in_data_reg_7,
	Add2,
	Add21,
	Add22,
	Add23,
	write_cp_data_77,
	write_cp_data_78,
	write_cp_data_75,
	write_cp_data_74,
	write_cp_data_76,
	WideNor0,
	nxt_out_eop,
	Equal14,
	src14_valid,
	src_valid,
	cp_ready1,
	in_data_reg_69,
	src_valid1,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_6,
	sink0_endofpacket,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	Selector3,
	Selector10,
	base_address_3,
	Selector4,
	Selector11,
	base_address_2,
	Selector5,
	Selector12,
	out_data_1,
	out_data_0,
	Selector6,
	Selector13,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARADDR_0;
input 	h2f_ARADDR_1;
input 	h2f_ARADDR_2;
input 	h2f_ARADDR_3;
input 	h2f_ARLEN_0;
output 	nxt_in_ready;
input 	in_ready_hold;
output 	stateST_COMP_TRANS;
output 	out_valid_reg1;
output 	in_narrow_reg1;
output 	in_byteen_reg_3;
output 	in_byteen_reg_2;
output 	in_byteen_reg_1;
output 	in_byteen_reg_0;
output 	in_data_reg_68;
input 	cp_ready;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready1;
input 	[128:0] sink0_data;
input 	Equal13;
input 	altera_reset_synchronizer_int_chain_out;
output 	in_data_reg_0;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
output 	in_data_reg_1;
output 	in_data_reg_2;
output 	in_data_reg_3;
output 	in_data_reg_4;
output 	in_data_reg_5;
output 	in_data_reg_6;
output 	in_data_reg_7;
input 	Add2;
input 	Add21;
input 	Add22;
input 	Add23;
input 	write_cp_data_77;
input 	write_cp_data_78;
input 	write_cp_data_75;
input 	write_cp_data_74;
input 	write_cp_data_76;
input 	WideNor0;
output 	nxt_out_eop;
input 	Equal14;
input 	src14_valid;
input 	src_valid;
input 	cp_ready1;
output 	in_data_reg_69;
input 	src_valid1;
output 	out_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_6;
input 	sink0_endofpacket;
output 	in_data_reg_105;
output 	in_data_reg_106;
output 	in_data_reg_107;
output 	in_data_reg_108;
output 	in_data_reg_109;
output 	in_data_reg_110;
output 	in_data_reg_111;
output 	in_data_reg_112;
output 	in_data_reg_113;
output 	in_data_reg_114;
output 	in_data_reg_115;
output 	in_data_reg_116;
input 	Selector3;
input 	Selector10;
input 	base_address_3;
input 	Selector4;
input 	Selector11;
input 	base_address_2;
input 	Selector5;
input 	Selector12;
input 	out_data_1;
input 	out_data_0;
input 	Selector6;
input 	Selector13;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \align_address_to_size|LessThan0~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt~0_combout ;
wire \Add4~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt[5]~1_combout ;
wire \nxt_uncomp_subburst_byte_cnt[4]~2_combout ;
wire \nxt_uncomp_subburst_byte_cnt[3]~3_combout ;
wire \nxt_uncomp_subburst_byte_cnt[2]~4_combout ;
wire \nxt_uncomp_subburst_byte_cnt[6]~5_combout ;
wire \WideOr0~combout ;
wire \in_valid~combout ;
wire \Selector0~0_combout ;
wire \load_next_out_cmd~combout ;
wire \state.ST_IDLE~q ;
wire \Selector2~0_combout ;
wire \Selector2~1_combout ;
wire \Selector2~2_combout ;
wire \state.ST_UNCOMP_TRANS~q ;
wire \Selector1~2_combout ;
wire \Selector1~0_combout ;
wire \Selector1~3_combout ;
wire \int_bytes_remaining_reg[5]~q ;
wire \d0_int_bytes_remaining[2]~4_combout ;
wire \d0_int_bytes_remaining[2]~5_combout ;
wire \int_bytes_remaining_reg[2]~q ;
wire \d0_int_bytes_remaining[3]~6_combout ;
wire \d0_int_bytes_remaining[3]~7_combout ;
wire \int_bytes_remaining_reg[3]~q ;
wire \Add1~1_combout ;
wire \d0_int_bytes_remaining[4]~8_combout ;
wire \int_bytes_remaining_reg[4]~q ;
wire \Add1~0_combout ;
wire \d0_int_bytes_remaining[5]~0_combout ;
wire \d0_int_bytes_remaining[5]~1_combout ;
wire \int_bytes_remaining_reg[6]~q ;
wire \d0_int_bytes_remaining[6]~2_combout ;
wire \d0_int_bytes_remaining[6]~3_combout ;
wire \Equal0~0_combout ;
wire \new_burst_reg~0_combout ;
wire \new_burst_reg~q ;
wire \Selector1~1_combout ;
wire \WideNor0~0_combout ;
wire \NON_PIPELINED_INPUTS.load_next_cmd~combout ;
wire \in_bytecount_reg_zero~q ;
wire \nxt_out_valid~0_combout ;
wire \LessThan0~0_combout ;
wire \Selector3~0_combout ;
wire \in_size_reg[0]~q ;
wire \in_size_reg[2]~q ;
wire \in_size_reg[1]~q ;
wire \ShiftLeft0~0_combout ;
wire \ShiftLeft0~1_combout ;
wire \int_byte_cnt_narrow_reg[3]~q ;
wire \ShiftLeft0~2_combout ;
wire \int_byte_cnt_narrow_reg[2]~q ;
wire \ShiftLeft0~3_combout ;
wire \ShiftLeft0~4_combout ;
wire \int_byte_cnt_narrow_reg[1]~q ;
wire \int_byte_cnt_narrow_reg[0]~q ;
wire \Add0~13_sumout ;
wire \d0_int_nxt_addr[0]~3_combout ;
wire \in_burstwrap_reg[0]~q ;
wire \nxt_addr[0]~0_combout ;
wire \int_nxt_addr_reg[0]~q ;
wire \d0_int_nxt_addr[0]~4_combout ;
wire \int_nxt_addr_reg_dly[0]~q ;
wire \Add0~14 ;
wire \Add0~9_sumout ;
wire \in_burstwrap_reg[1]~q ;
wire \nxt_addr[1]~4_combout ;
wire \int_nxt_addr_reg[1]~q ;
wire \d0_int_nxt_addr[1]~7_combout ;
wire \d0_int_nxt_addr[1]~2_combout ;
wire \int_nxt_addr_reg_dly[1]~q ;
wire \Add0~10 ;
wire \Add0~6 ;
wire \Add0~1_sumout ;
wire \in_burstwrap_reg[3]~q ;
wire \nxt_addr[3]~12_combout ;
wire \int_nxt_addr_reg[3]~q ;
wire \d0_int_nxt_addr[3]~5_combout ;
wire \d0_int_nxt_addr[3]~0_combout ;
wire \Add0~5_sumout ;
wire \in_burstwrap_reg[2]~q ;
wire \nxt_addr[2]~8_combout ;
wire \int_nxt_addr_reg[2]~q ;
wire \d0_int_nxt_addr[2]~6_combout ;
wire \d0_int_nxt_addr[2]~1_combout ;
wire \in_eop_reg~q ;


spw_babasu_altera_merlin_address_alignment_13 align_address_to_size(
	.new_burst_reg(\new_burst_reg~q ),
	.src_data_86(sink0_data[86]),
	.in_size_reg_0(\in_size_reg[0]~q ),
	.ShiftLeft0(\ShiftLeft0~3_combout ),
	.LessThan0(\align_address_to_size|LessThan0~0_combout ));

cyclonev_lcell_comb \nxt_in_ready~1 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!in_ready_hold),
	.datac(!out_valid_reg1),
	.datad(!cp_ready),
	.datae(!stateST_COMP_TRANS),
	.dataf(!\new_burst_reg~q ),
	.datag(!stateST_UNCOMP_WR_SUBBURST),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~1 .extended_lut = "on";
defparam \nxt_in_ready~1 .lut_mask = 64'h2020F0F02020F0FF;
defparam \nxt_in_ready~1 .shared_arith = "off";

dffeas \state.ST_COMP_TRANS (
	.clk(clk_clk),
	.d(\Selector1~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_COMP_TRANS),
	.prn(vcc));
defparam \state.ST_COMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_COMP_TRANS .power_up = "low";

dffeas out_valid_reg(
	.clk(clk_clk),
	.d(\nxt_out_valid~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_valid_reg1),
	.prn(vcc));
defparam out_valid_reg.is_wysiwyg = "true";
defparam out_valid_reg.power_up = "low";

dffeas in_narrow_reg(
	.clk(clk_clk),
	.d(\LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_narrow_reg1),
	.prn(vcc));
defparam in_narrow_reg.is_wysiwyg = "true";
defparam in_narrow_reg.power_up = "low";

dffeas \in_byteen_reg[3] (
	.clk(clk_clk),
	.d(sink0_data[35]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_3),
	.prn(vcc));
defparam \in_byteen_reg[3] .is_wysiwyg = "true";
defparam \in_byteen_reg[3] .power_up = "low";

dffeas \in_byteen_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[34]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_2),
	.prn(vcc));
defparam \in_byteen_reg[2] .is_wysiwyg = "true";
defparam \in_byteen_reg[2] .power_up = "low";

dffeas \in_byteen_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[33]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_1),
	.prn(vcc));
defparam \in_byteen_reg[1] .is_wysiwyg = "true";
defparam \in_byteen_reg[1] .power_up = "low";

dffeas \in_byteen_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[32]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_0),
	.prn(vcc));
defparam \in_byteen_reg[0] .is_wysiwyg = "true";
defparam \in_byteen_reg[0] .power_up = "low";

dffeas \in_data_reg[68] (
	.clk(clk_clk),
	.d(sink0_data[68]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_68),
	.prn(vcc));
defparam \in_data_reg[68] .is_wysiwyg = "true";
defparam \in_data_reg[68] .power_up = "low";

dffeas \state.ST_UNCOMP_WR_SUBBURST (
	.clk(clk_clk),
	.d(\Selector3~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_UNCOMP_WR_SUBBURST),
	.prn(vcc));
defparam \state.ST_UNCOMP_WR_SUBBURST .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_WR_SUBBURST .power_up = "low";

cyclonev_lcell_comb \nxt_in_ready~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!out_valid_reg1),
	.datac(!cp_ready),
	.datad(!\state.ST_UNCOMP_TRANS~q ),
	.datae(!stateST_UNCOMP_WR_SUBBURST),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~0 .extended_lut = "off";
defparam \nxt_in_ready~0 .lut_mask = 64'h008A8A8A008A8A8A;
defparam \nxt_in_ready~0 .shared_arith = "off";

dffeas \in_data_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[0]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_0),
	.prn(vcc));
defparam \in_data_reg[0] .is_wysiwyg = "true";
defparam \in_data_reg[0] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[3] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[3]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_3),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[3] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[2] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[2]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_2),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[2] .power_up = "low";

dffeas \in_data_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[1]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_1),
	.prn(vcc));
defparam \in_data_reg[1] .is_wysiwyg = "true";
defparam \in_data_reg[1] .power_up = "low";

dffeas \in_data_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[2]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_2),
	.prn(vcc));
defparam \in_data_reg[2] .is_wysiwyg = "true";
defparam \in_data_reg[2] .power_up = "low";

dffeas \in_data_reg[3] (
	.clk(clk_clk),
	.d(sink0_data[3]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_3),
	.prn(vcc));
defparam \in_data_reg[3] .is_wysiwyg = "true";
defparam \in_data_reg[3] .power_up = "low";

dffeas \in_data_reg[4] (
	.clk(clk_clk),
	.d(sink0_data[4]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_4),
	.prn(vcc));
defparam \in_data_reg[4] .is_wysiwyg = "true";
defparam \in_data_reg[4] .power_up = "low";

dffeas \in_data_reg[5] (
	.clk(clk_clk),
	.d(sink0_data[5]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_5),
	.prn(vcc));
defparam \in_data_reg[5] .is_wysiwyg = "true";
defparam \in_data_reg[5] .power_up = "low";

dffeas \in_data_reg[6] (
	.clk(clk_clk),
	.d(sink0_data[6]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_6),
	.prn(vcc));
defparam \in_data_reg[6] .is_wysiwyg = "true";
defparam \in_data_reg[6] .power_up = "low";

dffeas \in_data_reg[7] (
	.clk(clk_clk),
	.d(sink0_data[7]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_7),
	.prn(vcc));
defparam \in_data_reg[7] .is_wysiwyg = "true";
defparam \in_data_reg[7] .power_up = "low";

cyclonev_lcell_comb \nxt_out_eop~0 (
	.dataa(!\in_eop_reg~q ),
	.datab(!stateST_COMP_TRANS),
	.datac(!\new_burst_reg~q ),
	.datad(!cp_ready),
	.datae(!\in_bytecount_reg_zero~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_out_eop),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_eop~0 .extended_lut = "off";
defparam \nxt_out_eop~0 .lut_mask = 64'h4447774744477747;
defparam \nxt_out_eop~0 .shared_arith = "off";

dffeas \in_data_reg[69] (
	.clk(clk_clk),
	.d(sink0_data[69]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_69),
	.prn(vcc));
defparam \in_data_reg[69] .is_wysiwyg = "true";
defparam \in_data_reg[69] .power_up = "low";

dffeas \out_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[5] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[5]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_5),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[5] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[5] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[4] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[4]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_4),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[4] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[4] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[3] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[3]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_3),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[3] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[3] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[2]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[6] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[6]~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_6),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[6] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[6] .power_up = "low";

dffeas \in_data_reg[105] (
	.clk(clk_clk),
	.d(sink0_data[105]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_105),
	.prn(vcc));
defparam \in_data_reg[105] .is_wysiwyg = "true";
defparam \in_data_reg[105] .power_up = "low";

dffeas \in_data_reg[106] (
	.clk(clk_clk),
	.d(sink0_data[106]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_106),
	.prn(vcc));
defparam \in_data_reg[106] .is_wysiwyg = "true";
defparam \in_data_reg[106] .power_up = "low";

dffeas \in_data_reg[107] (
	.clk(clk_clk),
	.d(sink0_data[107]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_107),
	.prn(vcc));
defparam \in_data_reg[107] .is_wysiwyg = "true";
defparam \in_data_reg[107] .power_up = "low";

dffeas \in_data_reg[108] (
	.clk(clk_clk),
	.d(sink0_data[108]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_108),
	.prn(vcc));
defparam \in_data_reg[108] .is_wysiwyg = "true";
defparam \in_data_reg[108] .power_up = "low";

dffeas \in_data_reg[109] (
	.clk(clk_clk),
	.d(sink0_data[109]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_109),
	.prn(vcc));
defparam \in_data_reg[109] .is_wysiwyg = "true";
defparam \in_data_reg[109] .power_up = "low";

dffeas \in_data_reg[110] (
	.clk(clk_clk),
	.d(sink0_data[110]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_110),
	.prn(vcc));
defparam \in_data_reg[110] .is_wysiwyg = "true";
defparam \in_data_reg[110] .power_up = "low";

dffeas \in_data_reg[111] (
	.clk(clk_clk),
	.d(sink0_data[111]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_111),
	.prn(vcc));
defparam \in_data_reg[111] .is_wysiwyg = "true";
defparam \in_data_reg[111] .power_up = "low";

dffeas \in_data_reg[112] (
	.clk(clk_clk),
	.d(sink0_data[112]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_112),
	.prn(vcc));
defparam \in_data_reg[112] .is_wysiwyg = "true";
defparam \in_data_reg[112] .power_up = "low";

dffeas \in_data_reg[113] (
	.clk(clk_clk),
	.d(sink0_data[113]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_113),
	.prn(vcc));
defparam \in_data_reg[113] .is_wysiwyg = "true";
defparam \in_data_reg[113] .power_up = "low";

dffeas \in_data_reg[114] (
	.clk(clk_clk),
	.d(sink0_data[114]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_114),
	.prn(vcc));
defparam \in_data_reg[114] .is_wysiwyg = "true";
defparam \in_data_reg[114] .power_up = "low";

dffeas \in_data_reg[115] (
	.clk(clk_clk),
	.d(sink0_data[115]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_115),
	.prn(vcc));
defparam \in_data_reg[115] .is_wysiwyg = "true";
defparam \in_data_reg[115] .power_up = "low";

dffeas \in_data_reg[116] (
	.clk(clk_clk),
	.d(sink0_data[116]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_116),
	.prn(vcc));
defparam \in_data_reg[116] .is_wysiwyg = "true";
defparam \in_data_reg[116] .power_up = "low";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt~0 (
	.dataa(!out_valid_reg1),
	.datab(!cp_ready),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt~0 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt~0 .lut_mask = 64'h1111111111111111;
defparam \nxt_uncomp_subburst_byte_cnt~0 .shared_arith = "off";

cyclonev_lcell_comb \Add4~0 (
	.dataa(!out_uncomp_byte_cnt_reg_4),
	.datab(!out_uncomp_byte_cnt_reg_3),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add4~0 .extended_lut = "off";
defparam \Add4~0 .lut_mask = 64'h0800080008000800;
defparam \Add4~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[5]~1 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!\Add4~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[5]~1 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[5]~1 .lut_mask = 64'h0F4EA5E40F4EA5E4;
defparam \nxt_uncomp_subburst_byte_cnt[5]~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[4]~2 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!out_uncomp_byte_cnt_reg_3),
	.datae(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.dataf(!out_uncomp_byte_cnt_reg_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[4]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[4]~2 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[4]~2 .lut_mask = 64'h0F0FE44E0F0F4E4E;
defparam \nxt_uncomp_subburst_byte_cnt[4]~2 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[3]~3 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!out_uncomp_byte_cnt_reg_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[3]~3 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[3]~3 .lut_mask = 64'h0FE40F4E0FE40F4E;
defparam \nxt_uncomp_subburst_byte_cnt[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[2]~4 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[2]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[2]~4 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[2]~4 .lut_mask = 64'h0EF40EF40EF40EF4;
defparam \nxt_uncomp_subburst_byte_cnt[2]~4 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[6]~5 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!\Add4~0_combout ),
	.dataf(!out_uncomp_byte_cnt_reg_6),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[6]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[6]~5 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[6]~5 .lut_mask = 64'h0044A0E4FFEE5F4E;
defparam \nxt_uncomp_subburst_byte_cnt[6]~5 .shared_arith = "off";

cyclonev_lcell_comb WideOr0(
	.dataa(!\nxt_uncomp_subburst_byte_cnt[5]~1_combout ),
	.datab(!\nxt_uncomp_subburst_byte_cnt[4]~2_combout ),
	.datac(!\nxt_uncomp_subburst_byte_cnt[3]~3_combout ),
	.datad(!\nxt_uncomp_subburst_byte_cnt[2]~4_combout ),
	.datae(!\nxt_uncomp_subburst_byte_cnt[6]~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr0.extended_lut = "off";
defparam WideOr0.lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam WideOr0.shared_arith = "off";

cyclonev_lcell_comb in_valid(
	.dataa(!in_ready_hold),
	.datab(!Equal14),
	.datac(!Equal13),
	.datad(!sink0_data[68]),
	.datae(!src14_valid),
	.dataf(!src_valid),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\in_valid~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam in_valid.extended_lut = "off";
defparam in_valid.lut_mask = 64'h0000000155555555;
defparam in_valid.shared_arith = "off";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!sink0_data[69]),
	.datab(!nxt_out_eop),
	.datac(!sink0_data[68]),
	.datad(!\in_valid~combout ),
	.datae(!\state.ST_IDLE~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'h005FCCFF005FCCFF;
defparam \Selector0~0 .shared_arith = "off";

cyclonev_lcell_comb load_next_out_cmd(
	.dataa(!out_valid_reg1),
	.datab(!cp_ready),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\load_next_out_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam load_next_out_cmd.extended_lut = "off";
defparam load_next_out_cmd.lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam load_next_out_cmd.shared_arith = "off";

dffeas \state.ST_IDLE (
	.clk(clk_clk),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_IDLE~q ),
	.prn(vcc));
defparam \state.ST_IDLE .is_wysiwyg = "true";
defparam \state.ST_IDLE .power_up = "low";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!nxt_out_eop),
	.datac(!stateST_UNCOMP_WR_SUBBURST),
	.datad(!\state.ST_IDLE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'h00EC00EC00EC00EC;
defparam \Selector2~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~1 (
	.dataa(!in_ready_hold),
	.datab(!Equal14),
	.datac(!Equal13),
	.datad(!sink0_data[68]),
	.datae(!src14_valid),
	.dataf(!\Selector2~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~1 .extended_lut = "off";
defparam \Selector2~1 .lut_mask = 64'h0000000100000000;
defparam \Selector2~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~2 (
	.dataa(!\WideOr0~combout ),
	.datab(!\Selector2~1_combout ),
	.datac(!\in_valid~combout ),
	.datad(!nxt_out_eop),
	.datae(!\state.ST_UNCOMP_TRANS~q ),
	.dataf(!sink0_data[69]),
	.datag(!stateST_UNCOMP_WR_SUBBURST),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~2 .extended_lut = "on";
defparam \Selector2~2 .lut_mask = 64'h3B33BB3F0A00AA00;
defparam \Selector2~2 .shared_arith = "off";

dffeas \state.ST_UNCOMP_TRANS (
	.clk(clk_clk),
	.d(\Selector2~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_UNCOMP_TRANS~q ),
	.prn(vcc));
defparam \state.ST_UNCOMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_TRANS .power_up = "low";

cyclonev_lcell_comb \Selector1~2 (
	.dataa(!in_ready_hold),
	.datab(!stateST_COMP_TRANS),
	.datac(!nxt_out_eop),
	.datad(!sink0_data[68]),
	.datae(gnd),
	.dataf(!src_valid),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~2 .extended_lut = "off";
defparam \Selector1~2 .lut_mask = 64'h3030303031303130;
defparam \Selector1~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!nxt_out_eop),
	.datac(!\state.ST_UNCOMP_TRANS~q ),
	.datad(!stateST_UNCOMP_WR_SUBBURST),
	.datae(!\state.ST_IDLE~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'h0000A8880000A888;
defparam \Selector1~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~3 (
	.dataa(!in_ready_hold),
	.datab(!sink0_data[69]),
	.datac(!src_valid),
	.datad(!src_valid1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~3 .extended_lut = "off";
defparam \Selector1~3 .lut_mask = 64'h0111011101110111;
defparam \Selector1~3 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[5] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[5]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[5]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[5] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[5] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[2]~4 (
	.dataa(!h2f_ARLEN_0),
	.datab(!sink0_data[69]),
	.datac(!sink0_data[68]),
	.datad(!write_cp_data_74),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[2]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[2]~4 .extended_lut = "off";
defparam \d0_int_bytes_remaining[2]~4 .lut_mask = 64'h2F222F222F222F22;
defparam \d0_int_bytes_remaining[2]~4 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[2]~5 (
	.dataa(!\new_burst_reg~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\int_bytes_remaining_reg[2]~q ),
	.datad(!\d0_int_bytes_remaining[2]~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[2]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[2]~5 .extended_lut = "off";
defparam \d0_int_bytes_remaining[2]~5 .lut_mask = 64'h287D287D287D287D;
defparam \d0_int_bytes_remaining[2]~5 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[2] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[2]~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[2]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[2] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[3]~6 (
	.dataa(!sink0_data[69]),
	.datab(!sink0_data[68]),
	.datac(!write_cp_data_75),
	.datad(!Add2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[3]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[3]~6 .extended_lut = "off";
defparam \d0_int_bytes_remaining[3]~6 .lut_mask = 64'h0357035703570357;
defparam \d0_int_bytes_remaining[3]~6 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[3]~7 (
	.dataa(!\new_burst_reg~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\int_bytes_remaining_reg[2]~q ),
	.datad(!\int_bytes_remaining_reg[3]~q ),
	.datae(!\d0_int_bytes_remaining[3]~6_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[3]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[3]~7 .extended_lut = "off";
defparam \d0_int_bytes_remaining[3]~7 .lut_mask = 64'h208A75DF208A75DF;
defparam \d0_int_bytes_remaining[3]~7 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[3] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[3]~7_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[3]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[3] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[3] .power_up = "low";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!out_byte_cnt_reg_2),
	.datab(!\int_bytes_remaining_reg[2]~q ),
	.datac(!\int_bytes_remaining_reg[3]~q ),
	.datad(!\int_bytes_remaining_reg[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'hBF40BF40BF40BF40;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[4]~8 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!sink0_data[68]),
	.datad(!write_cp_data_76),
	.datae(!Add21),
	.dataf(!\Add1~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[4]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[4]~8 .extended_lut = "off";
defparam \d0_int_bytes_remaining[4]~8 .lut_mask = 64'hCCCFDDDF00031113;
defparam \d0_int_bytes_remaining[4]~8 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[4] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[4]~8_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[4]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[4] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[4] .power_up = "low";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!out_byte_cnt_reg_2),
	.datab(!\int_bytes_remaining_reg[2]~q ),
	.datac(!\int_bytes_remaining_reg[3]~q ),
	.datad(!\int_bytes_remaining_reg[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h4000400040004000;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[5]~0 (
	.dataa(!sink0_data[69]),
	.datab(!sink0_data[68]),
	.datac(!write_cp_data_77),
	.datad(!Add22),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[5]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[5]~0 .extended_lut = "off";
defparam \d0_int_bytes_remaining[5]~0 .lut_mask = 64'h0357035703570357;
defparam \d0_int_bytes_remaining[5]~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[5]~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\int_bytes_remaining_reg[5]~q ),
	.datac(!\Add1~0_combout ),
	.datad(!\d0_int_bytes_remaining[5]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[5]~1 .extended_lut = "off";
defparam \d0_int_bytes_remaining[5]~1 .lut_mask = 64'h287D287D287D287D;
defparam \d0_int_bytes_remaining[5]~1 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[6] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[6]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[6]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[6] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[6] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[6]~2 (
	.dataa(!sink0_data[69]),
	.datab(!sink0_data[68]),
	.datac(!write_cp_data_78),
	.datad(!Add23),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[6]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[6]~2 .extended_lut = "off";
defparam \d0_int_bytes_remaining[6]~2 .lut_mask = 64'h0357035703570357;
defparam \d0_int_bytes_remaining[6]~2 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[6]~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\int_bytes_remaining_reg[5]~q ),
	.datac(!\Add1~0_combout ),
	.datad(!\int_bytes_remaining_reg[6]~q ),
	.datae(!\d0_int_bytes_remaining[6]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[6]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[6]~3 .extended_lut = "off";
defparam \d0_int_bytes_remaining[6]~3 .lut_mask = 64'h08A25DF708A25DF7;
defparam \d0_int_bytes_remaining[6]~3 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!\d0_int_bytes_remaining[2]~5_combout ),
	.datab(!\d0_int_bytes_remaining[3]~7_combout ),
	.datac(!\d0_int_bytes_remaining[4]~8_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'h4040404040404040;
defparam \Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \new_burst_reg~0 (
	.dataa(!\Selector1~2_combout ),
	.datab(!\Selector1~0_combout ),
	.datac(!\Selector1~3_combout ),
	.datad(!\d0_int_bytes_remaining[5]~1_combout ),
	.datae(!\d0_int_bytes_remaining[6]~3_combout ),
	.dataf(!\Equal0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\new_burst_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \new_burst_reg~0 .extended_lut = "off";
defparam \new_burst_reg~0 .lut_mask = 64'hA2A2A2A2FFA2A2A2;
defparam \new_burst_reg~0 .shared_arith = "off";

dffeas new_burst_reg(
	.clk(clk_clk),
	.d(\new_burst_reg~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\new_burst_reg~q ),
	.prn(vcc));
defparam new_burst_reg.is_wysiwyg = "true";
defparam new_burst_reg.power_up = "low";

cyclonev_lcell_comb \Selector1~1 (
	.dataa(!sink0_data[69]),
	.datab(!stateST_COMP_TRANS),
	.datac(!nxt_out_eop),
	.datad(!sink0_data[68]),
	.datae(!\in_valid~combout ),
	.dataf(!\Selector1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~1 .extended_lut = "off";
defparam \Selector1~1 .lut_mask = 64'h3030777530303330;
defparam \Selector1~1 .shared_arith = "off";

cyclonev_lcell_comb \WideNor0~0 (
	.dataa(!sink0_data[69]),
	.datab(!sink0_data[68]),
	.datac(!WideNor0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideNor0~0 .extended_lut = "off";
defparam \WideNor0~0 .lut_mask = 64'h8A8A8A8A8A8A8A8A;
defparam \WideNor0~0 .shared_arith = "off";

cyclonev_lcell_comb \NON_PIPELINED_INPUTS.load_next_cmd (
	.dataa(!in_ready_hold),
	.datab(!nxt_in_ready1),
	.datac(!nxt_in_ready),
	.datad(!src_valid),
	.datae(!src_valid1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \NON_PIPELINED_INPUTS.load_next_cmd .extended_lut = "off";
defparam \NON_PIPELINED_INPUTS.load_next_cmd .lut_mask = 64'h0015151500151515;
defparam \NON_PIPELINED_INPUTS.load_next_cmd .shared_arith = "off";

dffeas in_bytecount_reg_zero(
	.clk(clk_clk),
	.d(\WideNor0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_bytecount_reg_zero~q ),
	.prn(vcc));
defparam in_bytecount_reg_zero.is_wysiwyg = "true";
defparam in_bytecount_reg_zero.power_up = "low";

cyclonev_lcell_comb \nxt_out_valid~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!\new_burst_reg~q ),
	.datac(!\in_bytecount_reg_zero~q ),
	.datad(!\in_valid~combout ),
	.datae(!cp_ready1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_valid~0 .extended_lut = "off";
defparam \nxt_out_valid~0 .lut_mask = 64'h50FF44FF50FF44FF;
defparam \nxt_out_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!sink0_data[87]),
	.datab(!sink0_data[88]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h8888888888888888;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~0 (
	.dataa(!nxt_out_eop),
	.datab(!\state.ST_UNCOMP_TRANS~q ),
	.datac(!stateST_UNCOMP_WR_SUBBURST),
	.datad(!\WideOr0~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'h002A002A002A002A;
defparam \Selector3~0 .shared_arith = "off";

dffeas \in_size_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[86]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[0]~q ),
	.prn(vcc));
defparam \in_size_reg[0] .is_wysiwyg = "true";
defparam \in_size_reg[0] .power_up = "low";

dffeas \in_size_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[88]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[2]~q ),
	.prn(vcc));
defparam \in_size_reg[2] .is_wysiwyg = "true";
defparam \in_size_reg[2] .power_up = "low";

dffeas \in_size_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[87]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[1]~q ),
	.prn(vcc));
defparam \in_size_reg[1] .is_wysiwyg = "true";
defparam \in_size_reg[1] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[87]),
	.datac(!sink0_data[88]),
	.datad(!\in_size_reg[2]~q ),
	.datae(!\in_size_reg[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~0 .extended_lut = "off";
defparam \ShiftLeft0~0 .lut_mask = 64'h1010BA101010BA10;
defparam \ShiftLeft0~0 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~1 .extended_lut = "off";
defparam \ShiftLeft0~1 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~1 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[3] (
	.clk(clk_clk),
	.d(\ShiftLeft0~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[3]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[3] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[3] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~2 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~2 .extended_lut = "off";
defparam \ShiftLeft0~2 .lut_mask = 64'h00E400E400E400E4;
defparam \ShiftLeft0~2 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[2] (
	.clk(clk_clk),
	.d(\ShiftLeft0~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[2]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[2] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[2] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[87]),
	.datac(!sink0_data[88]),
	.datad(!\in_size_reg[2]~q ),
	.datae(!\in_size_reg[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~3 .extended_lut = "off";
defparam \ShiftLeft0~3 .lut_mask = 64'hEA404040EA404040;
defparam \ShiftLeft0~3 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~4 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~4 .extended_lut = "off";
defparam \ShiftLeft0~4 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~4 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[1] (
	.clk(clk_clk),
	.d(\ShiftLeft0~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[1]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[1] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[1] .power_up = "low";

dffeas \int_byte_cnt_narrow_reg[0] (
	.clk(clk_clk),
	.d(\align_address_to_size|LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[0]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[0] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[0] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[0]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~3 (
	.dataa(!h2f_ARADDR_0),
	.datab(!sink0_data[69]),
	.datac(!sink0_data[68]),
	.datad(!out_data_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~3 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~3 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[0]~3 .shared_arith = "off";

dffeas \in_burstwrap_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[79]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[0]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[0] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[0] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[0]~0 (
	.dataa(!Selector13),
	.datab(!Selector6),
	.datac(!sink0_data[68]),
	.datad(!sink0_data[69]),
	.datae(!\new_burst_reg~q ),
	.dataf(!\d0_int_nxt_addr[0]~4_combout ),
	.datag(!\in_burstwrap_reg[0]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[0]~0 .extended_lut = "on";
defparam \nxt_addr[0]~0 .lut_mask = 64'h00000000F0F0FCA8;
defparam \nxt_addr[0]~0 .shared_arith = "off";

dffeas \int_nxt_addr_reg[0] (
	.clk(clk_clk),
	.d(\nxt_addr[0]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[0] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~4 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\Add0~13_sumout ),
	.datac(!\align_address_to_size|LessThan0~0_combout ),
	.datad(!\d0_int_nxt_addr[0]~3_combout ),
	.datae(!\int_nxt_addr_reg[0]~q ),
	.dataf(!\in_burstwrap_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~4 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~4 .lut_mask = 64'h0005AAAF2227AAAF;
defparam \d0_int_nxt_addr[0]~4 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[0] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[0]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[0] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[1]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[1]~q ),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \in_burstwrap_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[80]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[1]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[1] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[1] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[1]~4 (
	.dataa(!Selector12),
	.datab(!Selector5),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!\new_burst_reg~q ),
	.dataf(!\d0_int_nxt_addr[1]~2_combout ),
	.datag(!\in_burstwrap_reg[1]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[1]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[1]~4 .extended_lut = "on";
defparam \nxt_addr[1]~4 .lut_mask = 64'h00000000F0F0FAC8;
defparam \nxt_addr[1]~4 .shared_arith = "off";

dffeas \int_nxt_addr_reg[1] (
	.clk(clk_clk),
	.d(\nxt_addr[1]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[1] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~7 (
	.dataa(!h2f_ARADDR_1),
	.datab(!sink0_data[69]),
	.datac(!sink0_data[68]),
	.datad(!out_data_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~7 .extended_lut = "off";
defparam \d0_int_nxt_addr[1]~7 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[1]~7 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~2 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\Add0~9_sumout ),
	.datac(!\in_burstwrap_reg[1]~q ),
	.datad(!\int_nxt_addr_reg[1]~q ),
	.datae(!\ShiftLeft0~3_combout ),
	.dataf(!\d0_int_nxt_addr[1]~7_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~2 .extended_lut = "off";
defparam \d0_int_nxt_addr[1]~2 .lut_mask = 64'h02AA02AA02AA57FF;
defparam \d0_int_nxt_addr[1]~2 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[1] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[1]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[1] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_2),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[2]~q ),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[3]~q ),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

dffeas \in_burstwrap_reg[3] (
	.clk(clk_clk),
	.d(sink0_data[82]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[3]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[3] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[3] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[3]~12 (
	.dataa(!Selector10),
	.datab(!Selector3),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!\new_burst_reg~q ),
	.dataf(!\d0_int_nxt_addr[3]~0_combout ),
	.datag(!\in_burstwrap_reg[3]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[3]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[3]~12 .extended_lut = "on";
defparam \nxt_addr[3]~12 .lut_mask = 64'h00000000F0F0FAC8;
defparam \nxt_addr[3]~12 .shared_arith = "off";

dffeas \int_nxt_addr_reg[3] (
	.clk(clk_clk),
	.d(\nxt_addr[3]~12_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[3]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[3] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~5 (
	.dataa(!\Add0~1_sumout ),
	.datab(!\in_burstwrap_reg[3]~q ),
	.datac(!\int_nxt_addr_reg[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~5 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~5 .lut_mask = 64'hE0E0E0E0E0E0E0E0;
defparam \d0_int_nxt_addr[3]~5 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!h2f_ARADDR_3),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!base_address_3),
	.dataf(!\d0_int_nxt_addr[3]~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~0 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~0 .lut_mask = 64'hABABABFF01010155;
defparam \d0_int_nxt_addr[3]~0 .shared_arith = "off";

dffeas \in_burstwrap_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[81]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[2]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[2] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[2] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[2]~8 (
	.dataa(!Selector11),
	.datab(!Selector4),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!\new_burst_reg~q ),
	.dataf(!\d0_int_nxt_addr[2]~1_combout ),
	.datag(!\in_burstwrap_reg[2]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[2]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[2]~8 .extended_lut = "on";
defparam \nxt_addr[2]~8 .lut_mask = 64'h00000000F0F0FAC8;
defparam \nxt_addr[2]~8 .shared_arith = "off";

dffeas \int_nxt_addr_reg[2] (
	.clk(clk_clk),
	.d(\nxt_addr[2]~8_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[2]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~6 (
	.dataa(!\Add0~5_sumout ),
	.datab(!\in_burstwrap_reg[2]~q ),
	.datac(!\int_nxt_addr_reg[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~6 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~6 .lut_mask = 64'hE0E0E0E0E0E0E0E0;
defparam \d0_int_nxt_addr[2]~6 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!h2f_ARADDR_2),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!base_address_2),
	.dataf(!\d0_int_nxt_addr[2]~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~1 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~1 .lut_mask = 64'hABABABFF01010155;
defparam \d0_int_nxt_addr[2]~1 .shared_arith = "off";

dffeas in_eop_reg(
	.clk(clk_clk),
	.d(sink0_endofpacket),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_eop_reg~q ),
	.prn(vcc));
defparam in_eop_reg.is_wysiwyg = "true";
defparam in_eop_reg.power_up = "low";

endmodule

module spw_babasu_altera_merlin_address_alignment_13 (
	new_burst_reg,
	src_data_86,
	in_size_reg_0,
	ShiftLeft0,
	LessThan0)/* synthesis synthesis_greybox=0 */;
input 	new_burst_reg;
input 	src_data_86;
input 	in_size_reg_0;
input 	ShiftLeft0;
output 	LessThan0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!new_burst_reg),
	.datab(!src_data_86),
	.datac(!in_size_reg_0),
	.datad(!ShiftLeft0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan0),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h00E400E400E400E4;
defparam \LessThan0~0 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_burst_adapter_13 (
	h2f_ARADDR_0,
	h2f_ARADDR_1,
	h2f_ARADDR_2,
	h2f_ARADDR_3,
	h2f_ARBURST_0,
	h2f_ARBURST_1,
	h2f_ARID_0,
	h2f_ARID_1,
	h2f_ARID_2,
	h2f_ARID_3,
	h2f_ARID_4,
	h2f_ARID_5,
	h2f_ARID_6,
	h2f_ARID_7,
	h2f_ARID_8,
	h2f_ARID_9,
	h2f_ARID_10,
	h2f_ARID_11,
	h2f_ARLEN_0,
	Add5,
	Add51,
	Add52,
	in_ready_hold,
	saved_grant_1,
	stateST_COMP_TRANS,
	mem_used_1,
	in_data_reg_69,
	in_narrow_reg,
	cp_ready,
	cp_ready1,
	nxt_out_eop,
	out_valid_reg,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready,
	altera_reset_synchronizer_int_chain_out,
	Decoder1,
	Add2,
	Add21,
	Add22,
	Add23,
	nxt_in_ready1,
	src_valid,
	out_byte_cnt_reg_2,
	cp_ready2,
	out_uncomp_byte_cnt_reg_6,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	Selector10,
	Selector101,
	Add3,
	Add31,
	Selector11,
	Selector111,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	Add32,
	Selector12,
	src_payload,
	src_payload1,
	src_payload2,
	Selector13,
	nxt_out_burstwrap_1,
	nxt_addr_2,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARADDR_0;
input 	h2f_ARADDR_1;
input 	h2f_ARADDR_2;
input 	h2f_ARADDR_3;
input 	h2f_ARBURST_0;
input 	h2f_ARBURST_1;
input 	h2f_ARID_0;
input 	h2f_ARID_1;
input 	h2f_ARID_2;
input 	h2f_ARID_3;
input 	h2f_ARID_4;
input 	h2f_ARID_5;
input 	h2f_ARID_6;
input 	h2f_ARID_7;
input 	h2f_ARID_8;
input 	h2f_ARID_9;
input 	h2f_ARID_10;
input 	h2f_ARID_11;
input 	h2f_ARLEN_0;
input 	Add5;
input 	Add51;
input 	Add52;
input 	in_ready_hold;
input 	saved_grant_1;
output 	stateST_COMP_TRANS;
input 	mem_used_1;
output 	in_data_reg_69;
output 	in_narrow_reg;
input 	cp_ready;
input 	cp_ready1;
output 	nxt_out_eop;
output 	out_valid_reg;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready;
input 	altera_reset_synchronizer_int_chain_out;
input 	Decoder1;
input 	Add2;
input 	Add21;
input 	Add22;
input 	Add23;
output 	nxt_in_ready1;
input 	src_valid;
output 	out_byte_cnt_reg_2;
input 	cp_ready2;
output 	out_uncomp_byte_cnt_reg_6;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	in_data_reg_105;
output 	in_data_reg_106;
output 	in_data_reg_107;
output 	in_data_reg_108;
output 	in_data_reg_109;
output 	in_data_reg_110;
output 	in_data_reg_111;
output 	in_data_reg_112;
output 	in_data_reg_113;
output 	in_data_reg_114;
output 	in_data_reg_115;
output 	in_data_reg_116;
input 	Selector10;
input 	Selector101;
input 	Add3;
input 	Add31;
input 	Selector11;
input 	Selector111;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
input 	Add32;
input 	Selector12;
input 	src_payload;
input 	src_payload1;
input 	src_payload2;
input 	Selector13;
output 	nxt_out_burstwrap_1;
output 	nxt_addr_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



spw_babasu_altera_merlin_burst_adapter_13_1_13 \altera_merlin_burst_adapter_13_1.burst_adapter (
	.h2f_ARADDR_0(h2f_ARADDR_0),
	.h2f_ARADDR_1(h2f_ARADDR_1),
	.h2f_ARADDR_2(h2f_ARADDR_2),
	.h2f_ARADDR_3(h2f_ARADDR_3),
	.h2f_ARBURST_0(h2f_ARBURST_0),
	.h2f_ARBURST_1(h2f_ARBURST_1),
	.sink0_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,h2f_ARID_11,h2f_ARID_10,h2f_ARID_9,h2f_ARID_8,h2f_ARID_7,h2f_ARID_6,h2f_ARID_5,h2f_ARID_4,h2f_ARID_3,h2f_ARID_2,h2f_ARID_1,h2f_ARID_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_payload2,src_payload1,src_payload,gnd,gnd,gnd,
Selector101,Selector111,Selector12,Selector13,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,saved_grant_1,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.h2f_ARLEN_0(h2f_ARLEN_0),
	.Add5(Add5),
	.Add51(Add51),
	.Add52(Add52),
	.in_ready_hold(in_ready_hold),
	.stateST_COMP_TRANS(stateST_COMP_TRANS),
	.mem_used_1(mem_used_1),
	.in_data_reg_69(in_data_reg_69),
	.in_narrow_reg1(in_narrow_reg),
	.cp_ready(cp_ready),
	.cp_ready1(cp_ready1),
	.nxt_out_eop(nxt_out_eop),
	.out_valid_reg1(out_valid_reg),
	.stateST_UNCOMP_WR_SUBBURST(stateST_UNCOMP_WR_SUBBURST),
	.nxt_in_ready(nxt_in_ready),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.Decoder1(Decoder1),
	.Add2(Add2),
	.Add21(Add21),
	.Add22(Add22),
	.Add23(Add23),
	.nxt_in_ready1(nxt_in_ready1),
	.src_valid(src_valid),
	.out_byte_cnt_reg_2(out_byte_cnt_reg_2),
	.cp_ready2(cp_ready2),
	.out_uncomp_byte_cnt_reg_6(out_uncomp_byte_cnt_reg_6),
	.out_uncomp_byte_cnt_reg_5(out_uncomp_byte_cnt_reg_5),
	.out_uncomp_byte_cnt_reg_4(out_uncomp_byte_cnt_reg_4),
	.out_uncomp_byte_cnt_reg_3(out_uncomp_byte_cnt_reg_3),
	.out_uncomp_byte_cnt_reg_2(out_uncomp_byte_cnt_reg_2),
	.in_data_reg_105(in_data_reg_105),
	.in_data_reg_106(in_data_reg_106),
	.in_data_reg_107(in_data_reg_107),
	.in_data_reg_108(in_data_reg_108),
	.in_data_reg_109(in_data_reg_109),
	.in_data_reg_110(in_data_reg_110),
	.in_data_reg_111(in_data_reg_111),
	.in_data_reg_112(in_data_reg_112),
	.in_data_reg_113(in_data_reg_113),
	.in_data_reg_114(in_data_reg_114),
	.in_data_reg_115(in_data_reg_115),
	.in_data_reg_116(in_data_reg_116),
	.Selector10(Selector10),
	.Add3(Add3),
	.Add31(Add31),
	.Selector11(Selector11),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_3),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_2),
	.Add32(Add32),
	.nxt_out_burstwrap_1(nxt_out_burstwrap_1),
	.nxt_addr_2(nxt_addr_2),
	.clk_clk(clk_clk));

endmodule

module spw_babasu_altera_merlin_burst_adapter_13_1_13 (
	h2f_ARADDR_0,
	h2f_ARADDR_1,
	h2f_ARADDR_2,
	h2f_ARADDR_3,
	h2f_ARBURST_0,
	h2f_ARBURST_1,
	sink0_data,
	h2f_ARLEN_0,
	Add5,
	Add51,
	Add52,
	in_ready_hold,
	stateST_COMP_TRANS,
	mem_used_1,
	in_data_reg_69,
	in_narrow_reg1,
	cp_ready,
	cp_ready1,
	nxt_out_eop,
	out_valid_reg1,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready,
	altera_reset_synchronizer_int_chain_out,
	Decoder1,
	Add2,
	Add21,
	Add22,
	Add23,
	nxt_in_ready1,
	src_valid,
	out_byte_cnt_reg_2,
	cp_ready2,
	out_uncomp_byte_cnt_reg_6,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	Selector10,
	Add3,
	Add31,
	Selector11,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	Add32,
	nxt_out_burstwrap_1,
	nxt_addr_2,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARADDR_0;
input 	h2f_ARADDR_1;
input 	h2f_ARADDR_2;
input 	h2f_ARADDR_3;
input 	h2f_ARBURST_0;
input 	h2f_ARBURST_1;
input 	[128:0] sink0_data;
input 	h2f_ARLEN_0;
input 	Add5;
input 	Add51;
input 	Add52;
input 	in_ready_hold;
output 	stateST_COMP_TRANS;
input 	mem_used_1;
output 	in_data_reg_69;
output 	in_narrow_reg1;
input 	cp_ready;
input 	cp_ready1;
output 	nxt_out_eop;
output 	out_valid_reg1;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready;
input 	altera_reset_synchronizer_int_chain_out;
input 	Decoder1;
input 	Add2;
input 	Add21;
input 	Add22;
input 	Add23;
output 	nxt_in_ready1;
input 	src_valid;
output 	out_byte_cnt_reg_2;
input 	cp_ready2;
output 	out_uncomp_byte_cnt_reg_6;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	in_data_reg_105;
output 	in_data_reg_106;
output 	in_data_reg_107;
output 	in_data_reg_108;
output 	in_data_reg_109;
output 	in_data_reg_110;
output 	in_data_reg_111;
output 	in_data_reg_112;
output 	in_data_reg_113;
output 	in_data_reg_114;
output 	in_data_reg_115;
output 	in_data_reg_116;
input 	Selector10;
input 	Add3;
input 	Add31;
input 	Selector11;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
input 	Add32;
output 	nxt_out_burstwrap_1;
output 	nxt_addr_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \align_address_to_size|LessThan0~0_combout ;
wire \align_address_to_size|LessThan0~1_combout ;
wire \nxt_uncomp_subburst_byte_cnt~0_combout ;
wire \Add4~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt[6]~1_combout ;
wire \nxt_uncomp_subburst_byte_cnt[5]~2_combout ;
wire \nxt_uncomp_subburst_byte_cnt[4]~3_combout ;
wire \nxt_uncomp_subburst_byte_cnt[3]~4_combout ;
wire \nxt_uncomp_subburst_byte_cnt[2]~5_combout ;
wire \WideNor1~combout ;
wire \Selector2~1_combout ;
wire \load_next_out_cmd~combout ;
wire \state.ST_UNCOMP_TRANS~q ;
wire \Selector2~0_combout ;
wire \Selector0~0_combout ;
wire \state.ST_IDLE~q ;
wire \Selector1~0_combout ;
wire \Selector1~1_combout ;
wire \NON_PIPELINED_INPUTS.load_next_cmd~0_combout ;
wire \int_bytes_remaining_reg[4]~q ;
wire \d0_int_bytes_remaining[2]~3_combout ;
wire \int_bytes_remaining_reg[2]~q ;
wire \d0_int_bytes_remaining[3]~2_combout ;
wire \int_bytes_remaining_reg[3]~q ;
wire \Add1~0_combout ;
wire \d0_int_bytes_remaining[4]~0_combout ;
wire \int_bytes_remaining_reg[5]~q ;
wire \Add1~1_combout ;
wire \d0_int_bytes_remaining[5]~1_combout ;
wire \int_bytes_remaining_reg[6]~q ;
wire \d0_int_bytes_remaining[6]~4_combout ;
wire \new_burst_reg~0_combout ;
wire \new_burst_reg~q ;
wire \in_bytecount_reg_zero~0_combout ;
wire \in_bytecount_reg_zero~q ;
wire \nxt_out_valid~0_combout ;
wire \nxt_out_valid~1_combout ;
wire \Selector3~0_combout ;
wire \in_burstwrap_reg[3]~q ;
wire \nxt_addr[3]~0_combout ;
wire \nxt_addr[3]~combout ;
wire \int_nxt_addr_reg[3]~q ;
wire \in_size_reg[0]~q ;
wire \in_size_reg[1]~q ;
wire \in_size_reg[2]~q ;
wire \ShiftLeft0~0_combout ;
wire \ShiftLeft0~1_combout ;
wire \int_byte_cnt_narrow_reg[3]~q ;
wire \ShiftLeft0~2_combout ;
wire \int_byte_cnt_narrow_reg[2]~q ;
wire \in_burstwrap_reg[1]~q ;
wire \nxt_addr[1]~combout ;
wire \int_nxt_addr_reg[1]~q ;
wire \ShiftLeft0~3_combout ;
wire \int_byte_cnt_narrow_reg[1]~q ;
wire \int_byte_cnt_narrow_reg[0]~q ;
wire \Add0~13_sumout ;
wire \in_burstwrap_reg[0]~q ;
wire \nxt_addr[0]~combout ;
wire \int_nxt_addr_reg[0]~q ;
wire \d0_int_nxt_addr[0]~2_combout ;
wire \d0_int_nxt_addr[0]~3_combout ;
wire \int_nxt_addr_reg_dly[0]~q ;
wire \Add0~14 ;
wire \Add0~9_sumout ;
wire \d0_int_nxt_addr[1]~4_combout ;
wire \int_nxt_addr_reg_dly[1]~q ;
wire \Add0~10 ;
wire \Add0~6 ;
wire \Add0~1_sumout ;
wire \d0_int_nxt_addr[3]~0_combout ;
wire \in_burstwrap_reg[2]~q ;
wire \nxt_addr[2]~1_combout ;
wire \nxt_addr[2]~combout ;
wire \int_nxt_addr_reg[2]~q ;
wire \Add0~5_sumout ;
wire \d0_int_nxt_addr[2]~1_combout ;


spw_babasu_altera_merlin_address_alignment_14 align_address_to_size(
	.new_burst_reg(\new_burst_reg~q ),
	.src_payload(sink0_data[86]),
	.in_size_reg_0(\in_size_reg[0]~q ),
	.src_payload1(sink0_data[87]),
	.in_size_reg_1(\in_size_reg[1]~q ),
	.src_payload2(sink0_data[88]),
	.in_size_reg_2(\in_size_reg[2]~q ),
	.LessThan0(\align_address_to_size|LessThan0~0_combout ),
	.LessThan01(\align_address_to_size|LessThan0~1_combout ));

dffeas \state.ST_COMP_TRANS (
	.clk(clk_clk),
	.d(\Selector1~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_COMP_TRANS),
	.prn(vcc));
defparam \state.ST_COMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_COMP_TRANS .power_up = "low";

dffeas \in_data_reg[69] (
	.clk(clk_clk),
	.d(sink0_data[69]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_69),
	.prn(vcc));
defparam \in_data_reg[69] .is_wysiwyg = "true";
defparam \in_data_reg[69] .power_up = "low";

dffeas in_narrow_reg(
	.clk(clk_clk),
	.d(Decoder1),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_narrow_reg1),
	.prn(vcc));
defparam in_narrow_reg.is_wysiwyg = "true";
defparam in_narrow_reg.power_up = "low";

cyclonev_lcell_comb \nxt_out_eop~0 (
	.dataa(!in_data_reg_69),
	.datab(!stateST_COMP_TRANS),
	.datac(!\new_burst_reg~q ),
	.datad(!mem_used_1),
	.datae(!cp_ready),
	.dataf(!\in_bytecount_reg_zero~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_out_eop),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_eop~0 .extended_lut = "off";
defparam \nxt_out_eop~0 .lut_mask = 64'h4444474477774777;
defparam \nxt_out_eop~0 .shared_arith = "off";

dffeas out_valid_reg(
	.clk(clk_clk),
	.d(\nxt_out_valid~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_valid_reg1),
	.prn(vcc));
defparam out_valid_reg.is_wysiwyg = "true";
defparam out_valid_reg.power_up = "low";

dffeas \state.ST_UNCOMP_WR_SUBBURST (
	.clk(clk_clk),
	.d(\Selector3~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_UNCOMP_WR_SUBBURST),
	.prn(vcc));
defparam \state.ST_UNCOMP_WR_SUBBURST .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_WR_SUBBURST .power_up = "low";

cyclonev_lcell_comb \nxt_in_ready~0 (
	.dataa(!in_ready_hold),
	.datab(!stateST_COMP_TRANS),
	.datac(!mem_used_1),
	.datad(!cp_ready),
	.datae(!out_valid_reg1),
	.dataf(!\Selector2~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~0 .extended_lut = "off";
defparam \nxt_in_ready~0 .lut_mask = 64'h0000FF3F8888BBBB;
defparam \nxt_in_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_in_ready~1 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!cp_ready1),
	.datac(!nxt_out_eop),
	.datad(!nxt_in_ready),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~1 .extended_lut = "off";
defparam \nxt_in_ready~1 .lut_mask = 64'h00FE00FE00FE00FE;
defparam \nxt_in_ready~1 .shared_arith = "off";

dffeas \out_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[6] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[6]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_6),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[6] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[6] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[5] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[5]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_5),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[5] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[5] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[4] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[4]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_4),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[4] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[4] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[3] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[3]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_3),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[3] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[3] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[2]~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[2] .power_up = "low";

dffeas \in_data_reg[105] (
	.clk(clk_clk),
	.d(sink0_data[105]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_105),
	.prn(vcc));
defparam \in_data_reg[105] .is_wysiwyg = "true";
defparam \in_data_reg[105] .power_up = "low";

dffeas \in_data_reg[106] (
	.clk(clk_clk),
	.d(sink0_data[106]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_106),
	.prn(vcc));
defparam \in_data_reg[106] .is_wysiwyg = "true";
defparam \in_data_reg[106] .power_up = "low";

dffeas \in_data_reg[107] (
	.clk(clk_clk),
	.d(sink0_data[107]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_107),
	.prn(vcc));
defparam \in_data_reg[107] .is_wysiwyg = "true";
defparam \in_data_reg[107] .power_up = "low";

dffeas \in_data_reg[108] (
	.clk(clk_clk),
	.d(sink0_data[108]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_108),
	.prn(vcc));
defparam \in_data_reg[108] .is_wysiwyg = "true";
defparam \in_data_reg[108] .power_up = "low";

dffeas \in_data_reg[109] (
	.clk(clk_clk),
	.d(sink0_data[109]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_109),
	.prn(vcc));
defparam \in_data_reg[109] .is_wysiwyg = "true";
defparam \in_data_reg[109] .power_up = "low";

dffeas \in_data_reg[110] (
	.clk(clk_clk),
	.d(sink0_data[110]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_110),
	.prn(vcc));
defparam \in_data_reg[110] .is_wysiwyg = "true";
defparam \in_data_reg[110] .power_up = "low";

dffeas \in_data_reg[111] (
	.clk(clk_clk),
	.d(sink0_data[111]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_111),
	.prn(vcc));
defparam \in_data_reg[111] .is_wysiwyg = "true";
defparam \in_data_reg[111] .power_up = "low";

dffeas \in_data_reg[112] (
	.clk(clk_clk),
	.d(sink0_data[112]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_112),
	.prn(vcc));
defparam \in_data_reg[112] .is_wysiwyg = "true";
defparam \in_data_reg[112] .power_up = "low";

dffeas \in_data_reg[113] (
	.clk(clk_clk),
	.d(sink0_data[113]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_113),
	.prn(vcc));
defparam \in_data_reg[113] .is_wysiwyg = "true";
defparam \in_data_reg[113] .power_up = "low";

dffeas \in_data_reg[114] (
	.clk(clk_clk),
	.d(sink0_data[114]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_114),
	.prn(vcc));
defparam \in_data_reg[114] .is_wysiwyg = "true";
defparam \in_data_reg[114] .power_up = "low";

dffeas \in_data_reg[115] (
	.clk(clk_clk),
	.d(sink0_data[115]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_115),
	.prn(vcc));
defparam \in_data_reg[115] .is_wysiwyg = "true";
defparam \in_data_reg[115] .power_up = "low";

dffeas \in_data_reg[116] (
	.clk(clk_clk),
	.d(sink0_data[116]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_116),
	.prn(vcc));
defparam \in_data_reg[116] .is_wysiwyg = "true";
defparam \in_data_reg[116] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[3] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[3]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_3),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[3] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[2] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[2]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_2),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[2] .power_up = "low";

cyclonev_lcell_comb \nxt_out_burstwrap[1]~0 (
	.dataa(!h2f_ARBURST_0),
	.datab(!h2f_ARBURST_1),
	.datac(!Selector10),
	.datad(!Add32),
	.datae(!Add52),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_out_burstwrap_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_burstwrap[1]~0 .extended_lut = "off";
defparam \nxt_out_burstwrap[1]~0 .lut_mask = 64'h8A8802008A880200;
defparam \nxt_out_burstwrap[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_addr[2]~2 (
	.dataa(!Add3),
	.datab(!Add31),
	.datac(!Selector11),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_addr_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[2]~2 .extended_lut = "off";
defparam \nxt_addr[2]~2 .lut_mask = 64'h8080808080808080;
defparam \nxt_addr[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt~0 (
	.dataa(!cp_ready1),
	.datab(!out_valid_reg1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt~0 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt~0 .lut_mask = 64'h1111111111111111;
defparam \nxt_uncomp_subburst_byte_cnt~0 .shared_arith = "off";

cyclonev_lcell_comb \Add4~0 (
	.dataa(!out_uncomp_byte_cnt_reg_4),
	.datab(!out_uncomp_byte_cnt_reg_3),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add4~0 .extended_lut = "off";
defparam \Add4~0 .lut_mask = 64'h0800080008000800;
defparam \Add4~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[6]~1 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_6),
	.datad(!out_uncomp_byte_cnt_reg_5),
	.datae(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.dataf(!\Add4~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[6]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[6]~1 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[6]~1 .lut_mask = 64'h0F0F4E4EA50FE44E;
defparam \nxt_uncomp_subburst_byte_cnt[6]~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[5]~2 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!\Add4~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[5]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[5]~2 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[5]~2 .lut_mask = 64'h0F4EA5E40F4EA5E4;
defparam \nxt_uncomp_subburst_byte_cnt[5]~2 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[4]~3 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!out_uncomp_byte_cnt_reg_3),
	.datae(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.dataf(!out_uncomp_byte_cnt_reg_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[4]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[4]~3 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[4]~3 .lut_mask = 64'h0F0FE44E0F0F4E4E;
defparam \nxt_uncomp_subburst_byte_cnt[4]~3 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[3]~4 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!out_uncomp_byte_cnt_reg_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[3]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[3]~4 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[3]~4 .lut_mask = 64'h0FE40F4E0FE40F4E;
defparam \nxt_uncomp_subburst_byte_cnt[3]~4 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[2]~5 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[2]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[2]~5 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[2]~5 .lut_mask = 64'h0EF40EF40EF40EF4;
defparam \nxt_uncomp_subburst_byte_cnt[2]~5 .shared_arith = "off";

cyclonev_lcell_comb WideNor1(
	.dataa(!\nxt_uncomp_subburst_byte_cnt[6]~1_combout ),
	.datab(!\nxt_uncomp_subburst_byte_cnt[5]~2_combout ),
	.datac(!\nxt_uncomp_subburst_byte_cnt[4]~3_combout ),
	.datad(!\nxt_uncomp_subburst_byte_cnt[3]~4_combout ),
	.datae(!\nxt_uncomp_subburst_byte_cnt[2]~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideNor1.extended_lut = "off";
defparam WideNor1.lut_mask = 64'h8000000080000000;
defparam WideNor1.shared_arith = "off";

cyclonev_lcell_comb \Selector2~1 (
	.dataa(!nxt_out_eop),
	.datab(!\Selector2~0_combout ),
	.datac(!\WideNor1~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~1 .extended_lut = "off";
defparam \Selector2~1 .lut_mask = 64'h0808080808080808;
defparam \Selector2~1 .shared_arith = "off";

cyclonev_lcell_comb load_next_out_cmd(
	.dataa(!mem_used_1),
	.datab(!cp_ready),
	.datac(!out_valid_reg1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\load_next_out_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam load_next_out_cmd.extended_lut = "off";
defparam load_next_out_cmd.lut_mask = 64'hF2F2F2F2F2F2F2F2;
defparam load_next_out_cmd.shared_arith = "off";

dffeas \state.ST_UNCOMP_TRANS (
	.clk(clk_clk),
	.d(\Selector2~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_UNCOMP_TRANS~q ),
	.prn(vcc));
defparam \state.ST_UNCOMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_TRANS .power_up = "low";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'h8888888888888888;
defparam \Selector2~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!in_ready_hold),
	.datab(!nxt_out_eop),
	.datac(!src_valid),
	.datad(!\state.ST_IDLE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'h05CD05CD05CD05CD;
defparam \Selector0~0 .shared_arith = "off";

dffeas \state.ST_IDLE (
	.clk(clk_clk),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_IDLE~q ),
	.prn(vcc));
defparam \state.ST_IDLE .is_wysiwyg = "true";
defparam \state.ST_IDLE .power_up = "low";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!sink0_data[69]),
	.datab(!nxt_out_eop),
	.datac(!\Selector2~0_combout ),
	.datad(!\state.ST_IDLE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'h5510551055105510;
defparam \Selector1~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~1 (
	.dataa(!in_ready_hold),
	.datab(!stateST_COMP_TRANS),
	.datac(!nxt_out_eop),
	.datad(!src_valid),
	.datae(!\Selector1~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~1 .extended_lut = "off";
defparam \Selector1~1 .lut_mask = 64'h3031307530313075;
defparam \Selector1~1 .shared_arith = "off";

cyclonev_lcell_comb \NON_PIPELINED_INPUTS.load_next_cmd~0 (
	.dataa(!in_ready_hold),
	.datab(!nxt_in_ready1),
	.datac(!src_valid),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \NON_PIPELINED_INPUTS.load_next_cmd~0 .extended_lut = "off";
defparam \NON_PIPELINED_INPUTS.load_next_cmd~0 .lut_mask = 64'h0404040404040404;
defparam \NON_PIPELINED_INPUTS.load_next_cmd~0 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[4] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[4]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[4]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[4] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[4] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[2]~3 (
	.dataa(!h2f_ARLEN_0),
	.datab(!sink0_data[69]),
	.datac(!\new_burst_reg~q ),
	.datad(!out_byte_cnt_reg_2),
	.datae(!\int_bytes_remaining_reg[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[2]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[2]~3 .extended_lut = "off";
defparam \d0_int_bytes_remaining[2]~3 .lut_mask = 64'h02F2F20202F2F202;
defparam \d0_int_bytes_remaining[2]~3 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[2] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[2]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[2]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[2] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[3]~2 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!Add2),
	.datad(!\int_bytes_remaining_reg[3]~q ),
	.datae(!out_byte_cnt_reg_2),
	.dataf(!\int_bytes_remaining_reg[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[3]~2 .extended_lut = "off";
defparam \d0_int_bytes_remaining[3]~2 .lut_mask = 64'h01CDCD0101CD01CD;
defparam \d0_int_bytes_remaining[3]~2 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[3] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[3]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[3]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[3] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[3] .power_up = "low";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!\int_bytes_remaining_reg[4]~q ),
	.datab(!\int_bytes_remaining_reg[3]~q ),
	.datac(!out_byte_cnt_reg_2),
	.datad(!\int_bytes_remaining_reg[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'hA6AAA6AAA6AAA6AA;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[4]~0 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!Add21),
	.datad(!\Add1~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[4]~0 .extended_lut = "off";
defparam \d0_int_bytes_remaining[4]~0 .lut_mask = 64'hCD01CD01CD01CD01;
defparam \d0_int_bytes_remaining[4]~0 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[5] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[5]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[5]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[5] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[5] .power_up = "low";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!\int_bytes_remaining_reg[4]~q ),
	.datab(!\int_bytes_remaining_reg[3]~q ),
	.datac(!out_byte_cnt_reg_2),
	.datad(!\int_bytes_remaining_reg[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h0800080008000800;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[5]~1 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!Add22),
	.datad(!\int_bytes_remaining_reg[5]~q ),
	.datae(!\Add1~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[5]~1 .extended_lut = "off";
defparam \d0_int_bytes_remaining[5]~1 .lut_mask = 64'h01CDCD0101CDCD01;
defparam \d0_int_bytes_remaining[5]~1 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[6] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[6]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[6]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[6] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[6] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[6]~4 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!Add23),
	.datad(!\int_bytes_remaining_reg[5]~q ),
	.datae(!\Add1~1_combout ),
	.dataf(!\int_bytes_remaining_reg[6]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[6]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[6]~4 .extended_lut = "off";
defparam \d0_int_bytes_remaining[6]~4 .lut_mask = 64'h0101CD01CDCD01CD;
defparam \d0_int_bytes_remaining[6]~4 .shared_arith = "off";

cyclonev_lcell_comb \new_burst_reg~0 (
	.dataa(!\Selector1~1_combout ),
	.datab(!\d0_int_bytes_remaining[4]~0_combout ),
	.datac(!\d0_int_bytes_remaining[5]~1_combout ),
	.datad(!\d0_int_bytes_remaining[3]~2_combout ),
	.datae(!\d0_int_bytes_remaining[2]~3_combout ),
	.dataf(!\d0_int_bytes_remaining[6]~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\new_burst_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \new_burst_reg~0 .extended_lut = "off";
defparam \new_burst_reg~0 .lut_mask = 64'hAAAAEAAAAAAAAAAA;
defparam \new_burst_reg~0 .shared_arith = "off";

dffeas new_burst_reg(
	.clk(clk_clk),
	.d(\new_burst_reg~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\new_burst_reg~q ),
	.prn(vcc));
defparam new_burst_reg.is_wysiwyg = "true";
defparam new_burst_reg.power_up = "low";

cyclonev_lcell_comb \in_bytecount_reg_zero~0 (
	.dataa(!sink0_data[69]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\in_bytecount_reg_zero~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \in_bytecount_reg_zero~0 .extended_lut = "off";
defparam \in_bytecount_reg_zero~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \in_bytecount_reg_zero~0 .shared_arith = "off";

dffeas in_bytecount_reg_zero(
	.clk(clk_clk),
	.d(\in_bytecount_reg_zero~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_bytecount_reg_zero~q ),
	.prn(vcc));
defparam in_bytecount_reg_zero.is_wysiwyg = "true";
defparam in_bytecount_reg_zero.power_up = "low";

cyclonev_lcell_comb \nxt_out_valid~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!mem_used_1),
	.datac(!\in_bytecount_reg_zero~q ),
	.datad(!cp_ready2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_valid~0 .extended_lut = "off";
defparam \nxt_out_valid~0 .lut_mask = 64'hF0B8F0B8F0B8F0B8;
defparam \nxt_out_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_out_valid~1 (
	.dataa(!in_ready_hold),
	.datab(!stateST_COMP_TRANS),
	.datac(!src_valid),
	.datad(!\nxt_out_valid~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_valid~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_valid~1 .extended_lut = "off";
defparam \nxt_out_valid~1 .lut_mask = 64'h0537053705370537;
defparam \nxt_out_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~0 (
	.dataa(!nxt_out_eop),
	.datab(!\Selector2~0_combout ),
	.datac(!\WideNor1~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'h8080808080808080;
defparam \Selector3~0 .shared_arith = "off";

dffeas \in_burstwrap_reg[3] (
	.clk(clk_clk),
	.d(sink0_data[82]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_burstwrap_reg[3]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[3] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[3] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[3]~0 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!\in_burstwrap_reg[3]~q ),
	.datad(!\d0_int_nxt_addr[3]~0_combout ),
	.datae(!h2f_ARBURST_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[3]~0 .extended_lut = "off";
defparam \nxt_addr[3]~0 .lut_mask = 64'h00F300E200F300E2;
defparam \nxt_addr[3]~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_addr[3] (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!h2f_ARBURST_1),
	.datad(!Add5),
	.datae(!Selector10),
	.dataf(!\nxt_addr[3]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[3] .extended_lut = "off";
defparam \nxt_addr[3] .lut_mask = 64'h00000000FEEEFFEF;
defparam \nxt_addr[3] .shared_arith = "off";

dffeas \int_nxt_addr_reg[3] (
	.clk(clk_clk),
	.d(\nxt_addr[3]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[3]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[3] .power_up = "low";

dffeas \in_size_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[86]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_size_reg[0]~q ),
	.prn(vcc));
defparam \in_size_reg[0] .is_wysiwyg = "true";
defparam \in_size_reg[0] .power_up = "low";

dffeas \in_size_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[87]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_size_reg[1]~q ),
	.prn(vcc));
defparam \in_size_reg[1] .is_wysiwyg = "true";
defparam \in_size_reg[1] .power_up = "low";

dffeas \in_size_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[88]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_size_reg[2]~q ),
	.prn(vcc));
defparam \in_size_reg[2] .is_wysiwyg = "true";
defparam \in_size_reg[2] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[87]),
	.datac(!\in_size_reg[1]~q ),
	.datad(!sink0_data[88]),
	.datae(!\in_size_reg[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~0 .extended_lut = "off";
defparam \ShiftLeft0~0 .lut_mask = 64'h1B0A11001B0A1100;
defparam \ShiftLeft0~0 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~1 .extended_lut = "off";
defparam \ShiftLeft0~1 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~1 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[3] (
	.clk(clk_clk),
	.d(\ShiftLeft0~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[3]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[3] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[3] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~2 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~2 .extended_lut = "off";
defparam \ShiftLeft0~2 .lut_mask = 64'h00E400E400E400E4;
defparam \ShiftLeft0~2 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[2] (
	.clk(clk_clk),
	.d(\ShiftLeft0~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[2]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[2] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[2] .power_up = "low";

dffeas \in_burstwrap_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[80]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_burstwrap_reg[1]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[1] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[1] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[1] (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!\in_burstwrap_reg[1]~q ),
	.datad(!\d0_int_nxt_addr[1]~4_combout ),
	.datae(!nxt_out_burstwrap_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[1] .extended_lut = "off";
defparam \nxt_addr[1] .lut_mask = 64'h00E200F300E200F3;
defparam \nxt_addr[1] .shared_arith = "off";

dffeas \int_nxt_addr_reg[1] (
	.clk(clk_clk),
	.d(\nxt_addr[1]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[1] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\align_address_to_size|LessThan0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~3 .extended_lut = "off";
defparam \ShiftLeft0~3 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~3 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[1] (
	.clk(clk_clk),
	.d(\ShiftLeft0~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[1]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[1] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[1] .power_up = "low";

dffeas \int_byte_cnt_narrow_reg[0] (
	.clk(clk_clk),
	.d(\align_address_to_size|LessThan0~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[0]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[0] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[0] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[0]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \in_burstwrap_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[79]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_burstwrap_reg[0]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[0] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[0] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[0] (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!sink0_data[79]),
	.datad(!\in_burstwrap_reg[0]~q ),
	.datae(!\d0_int_nxt_addr[0]~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[0] .extended_lut = "off";
defparam \nxt_addr[0] .lut_mask = 64'h0000FE320000FE32;
defparam \nxt_addr[0] .shared_arith = "off";

dffeas \int_nxt_addr_reg[0] (
	.clk(clk_clk),
	.d(\nxt_addr[0]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[0] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~2 (
	.dataa(!\Add0~13_sumout ),
	.datab(!\int_nxt_addr_reg[0]~q ),
	.datac(!\in_burstwrap_reg[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~2 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~2 .lut_mask = 64'hC8C8C8C8C8C8C8C8;
defparam \d0_int_nxt_addr[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~3 (
	.dataa(!h2f_ARADDR_0),
	.datab(!sink0_data[69]),
	.datac(!\new_burst_reg~q ),
	.datad(!\align_address_to_size|LessThan0~1_combout ),
	.datae(!\d0_int_nxt_addr[0]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~3 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~3 .lut_mask = 64'hF0F10001F0F10001;
defparam \d0_int_nxt_addr[0]~3 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[0] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[0]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[0] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[1]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[1]~q ),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~4 (
	.dataa(!\int_nxt_addr_reg[1]~q ),
	.datab(!\Add0~9_sumout ),
	.datac(!sink0_data[69]),
	.datad(!Decoder1),
	.datae(!\new_burst_reg~q ),
	.dataf(!h2f_ARADDR_1),
	.datag(!\in_burstwrap_reg[1]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~4 .extended_lut = "on";
defparam \d0_int_nxt_addr[1]~4 .lut_mask = 64'h575700005757000F;
defparam \d0_int_nxt_addr[1]~4 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[1] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[1]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[1] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_2),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[2]~q ),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[3]~q ),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~0 (
	.dataa(!h2f_ARADDR_3),
	.datab(!sink0_data[69]),
	.datac(!\new_burst_reg~q ),
	.datad(!\int_nxt_addr_reg[3]~q ),
	.datae(!\in_burstwrap_reg[3]~q ),
	.dataf(!\Add0~1_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~0 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~0 .lut_mask = 64'h01F101F101F1F1F1;
defparam \d0_int_nxt_addr[3]~0 .shared_arith = "off";

dffeas \in_burstwrap_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[81]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_burstwrap_reg[2]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[2] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[2] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[2]~1 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!\in_burstwrap_reg[2]~q ),
	.datad(!\d0_int_nxt_addr[2]~1_combout ),
	.datae(!h2f_ARBURST_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[2]~1 .extended_lut = "off";
defparam \nxt_addr[2]~1 .lut_mask = 64'h00F300E200F300E2;
defparam \nxt_addr[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_addr[2] (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!h2f_ARBURST_1),
	.datad(!Add51),
	.datae(!\nxt_addr[2]~1_combout ),
	.dataf(!nxt_addr_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[2] .extended_lut = "off";
defparam \nxt_addr[2] .lut_mask = 64'h0000FEEE0000FFEF;
defparam \nxt_addr[2] .shared_arith = "off";

dffeas \int_nxt_addr_reg[2] (
	.clk(clk_clk),
	.d(\nxt_addr[2]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[2]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~1 (
	.dataa(!h2f_ARADDR_2),
	.datab(!sink0_data[69]),
	.datac(!\new_burst_reg~q ),
	.datad(!\int_nxt_addr_reg[2]~q ),
	.datae(!\in_burstwrap_reg[2]~q ),
	.dataf(!\Add0~5_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~1 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~1 .lut_mask = 64'h01F101F101F1F1F1;
defparam \d0_int_nxt_addr[2]~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_address_alignment_14 (
	new_burst_reg,
	src_payload,
	in_size_reg_0,
	src_payload1,
	in_size_reg_1,
	src_payload2,
	in_size_reg_2,
	LessThan0,
	LessThan01)/* synthesis synthesis_greybox=0 */;
input 	new_burst_reg;
input 	src_payload;
input 	in_size_reg_0;
input 	src_payload1;
input 	in_size_reg_1;
input 	src_payload2;
input 	in_size_reg_2;
output 	LessThan0;
output 	LessThan01;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!new_burst_reg),
	.datab(!src_payload1),
	.datac(!in_size_reg_1),
	.datad(!src_payload2),
	.datae(!in_size_reg_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan0),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'hE4A04400E4A04400;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~1 (
	.dataa(!new_burst_reg),
	.datab(!src_payload),
	.datac(!in_size_reg_0),
	.datad(!LessThan0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan01),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~1 .extended_lut = "off";
defparam \LessThan0~1 .lut_mask = 64'h00E400E400E400E4;
defparam \LessThan0~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_burst_adapter_14 (
	h2f_ARADDR_0,
	h2f_ARADDR_1,
	h2f_ARADDR_2,
	h2f_ARADDR_3,
	h2f_ARLEN_0,
	nxt_in_ready,
	in_ready_hold,
	stateST_COMP_TRANS,
	out_valid_reg,
	in_narrow_reg,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	in_data_reg_68,
	cp_ready,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready1,
	saved_grant_1,
	Equal15,
	saved_grant_0,
	altera_reset_synchronizer_int_chain_out,
	in_data_reg_0,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	in_data_reg_1,
	in_data_reg_2,
	in_data_reg_3,
	in_data_reg_4,
	in_data_reg_5,
	in_data_reg_6,
	Add2,
	Add21,
	Add22,
	Add23,
	write_cp_data_77,
	write_cp_data_78,
	write_cp_data_75,
	write_cp_data_74,
	write_cp_data_76,
	WideNor0,
	nxt_out_eop,
	Equal151,
	src15_valid,
	src_valid,
	cp_ready1,
	in_data_reg_69,
	src_data_87,
	src_data_88,
	src_valid1,
	src_data_35,
	src_data_34,
	src_data_33,
	src_data_32,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_6,
	src_payload_0,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	Selector3,
	Selector10,
	base_address_3,
	Selector4,
	Selector11,
	base_address_2,
	src_payload,
	src_data_82,
	src_data_81,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_data_105,
	src_data_106,
	src_data_107,
	src_data_108,
	src_data_109,
	src_data_110,
	src_data_111,
	src_data_112,
	src_data_113,
	src_data_114,
	src_data_115,
	src_data_116,
	src_data_86,
	Selector5,
	Selector12,
	out_data_1,
	src_data_80,
	out_data_0,
	Selector6,
	Selector13,
	src_data_79,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARADDR_0;
input 	h2f_ARADDR_1;
input 	h2f_ARADDR_2;
input 	h2f_ARADDR_3;
input 	h2f_ARLEN_0;
output 	nxt_in_ready;
input 	in_ready_hold;
output 	stateST_COMP_TRANS;
output 	out_valid_reg;
output 	in_narrow_reg;
output 	in_byteen_reg_3;
output 	in_byteen_reg_2;
output 	in_byteen_reg_1;
output 	in_byteen_reg_0;
output 	in_data_reg_68;
input 	cp_ready;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready1;
input 	saved_grant_1;
input 	Equal15;
input 	saved_grant_0;
input 	altera_reset_synchronizer_int_chain_out;
output 	in_data_reg_0;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
output 	in_data_reg_1;
output 	in_data_reg_2;
output 	in_data_reg_3;
output 	in_data_reg_4;
output 	in_data_reg_5;
output 	in_data_reg_6;
input 	Add2;
input 	Add21;
input 	Add22;
input 	Add23;
input 	write_cp_data_77;
input 	write_cp_data_78;
input 	write_cp_data_75;
input 	write_cp_data_74;
input 	write_cp_data_76;
input 	WideNor0;
output 	nxt_out_eop;
input 	Equal151;
input 	src15_valid;
input 	src_valid;
input 	cp_ready1;
output 	in_data_reg_69;
input 	src_data_87;
input 	src_data_88;
input 	src_valid1;
input 	src_data_35;
input 	src_data_34;
input 	src_data_33;
input 	src_data_32;
output 	out_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_6;
input 	src_payload_0;
output 	in_data_reg_105;
output 	in_data_reg_106;
output 	in_data_reg_107;
output 	in_data_reg_108;
output 	in_data_reg_109;
output 	in_data_reg_110;
output 	in_data_reg_111;
output 	in_data_reg_112;
output 	in_data_reg_113;
output 	in_data_reg_114;
output 	in_data_reg_115;
output 	in_data_reg_116;
input 	Selector3;
input 	Selector10;
input 	base_address_3;
input 	Selector4;
input 	Selector11;
input 	base_address_2;
input 	src_payload;
input 	src_data_82;
input 	src_data_81;
input 	src_payload1;
input 	src_payload2;
input 	src_payload3;
input 	src_payload4;
input 	src_payload5;
input 	src_payload6;
input 	src_data_105;
input 	src_data_106;
input 	src_data_107;
input 	src_data_108;
input 	src_data_109;
input 	src_data_110;
input 	src_data_111;
input 	src_data_112;
input 	src_data_113;
input 	src_data_114;
input 	src_data_115;
input 	src_data_116;
input 	src_data_86;
input 	Selector5;
input 	Selector12;
input 	out_data_1;
input 	src_data_80;
input 	out_data_0;
input 	Selector6;
input 	Selector13;
input 	src_data_79;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



spw_babasu_altera_merlin_burst_adapter_13_1_14 \altera_merlin_burst_adapter_13_1.burst_adapter (
	.h2f_ARADDR_0(h2f_ARADDR_0),
	.h2f_ARADDR_1(h2f_ARADDR_1),
	.h2f_ARADDR_2(h2f_ARADDR_2),
	.h2f_ARADDR_3(h2f_ARADDR_3),
	.h2f_ARLEN_0(h2f_ARLEN_0),
	.nxt_in_ready(nxt_in_ready),
	.in_ready_hold(in_ready_hold),
	.stateST_COMP_TRANS(stateST_COMP_TRANS),
	.out_valid_reg1(out_valid_reg),
	.in_narrow_reg1(in_narrow_reg),
	.in_byteen_reg_3(in_byteen_reg_3),
	.in_byteen_reg_2(in_byteen_reg_2),
	.in_byteen_reg_1(in_byteen_reg_1),
	.in_byteen_reg_0(in_byteen_reg_0),
	.in_data_reg_68(in_data_reg_68),
	.cp_ready(cp_ready),
	.stateST_UNCOMP_WR_SUBBURST(stateST_UNCOMP_WR_SUBBURST),
	.nxt_in_ready1(nxt_in_ready1),
	.sink0_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_116,src_data_115,src_data_114,src_data_113,src_data_112,src_data_111,src_data_110,src_data_109,src_data_108,src_data_107,src_data_106,src_data_105,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_88,src_data_87,
src_data_86,gnd,gnd,gnd,src_data_82,src_data_81,src_data_80,src_data_79,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,saved_grant_1,saved_grant_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_35,src_data_34,src_data_33,
src_data_32,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_payload6,src_payload5,src_payload4,src_payload3,src_payload2,src_payload1,src_payload}),
	.Equal15(Equal15),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.in_data_reg_0(in_data_reg_0),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_3),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_2),
	.in_data_reg_1(in_data_reg_1),
	.in_data_reg_2(in_data_reg_2),
	.in_data_reg_3(in_data_reg_3),
	.in_data_reg_4(in_data_reg_4),
	.in_data_reg_5(in_data_reg_5),
	.in_data_reg_6(in_data_reg_6),
	.Add2(Add2),
	.Add21(Add21),
	.Add22(Add22),
	.Add23(Add23),
	.write_cp_data_77(write_cp_data_77),
	.write_cp_data_78(write_cp_data_78),
	.write_cp_data_75(write_cp_data_75),
	.write_cp_data_74(write_cp_data_74),
	.write_cp_data_76(write_cp_data_76),
	.WideNor0(WideNor0),
	.nxt_out_eop(nxt_out_eop),
	.Equal151(Equal151),
	.src15_valid(src15_valid),
	.src_valid(src_valid),
	.cp_ready1(cp_ready1),
	.in_data_reg_69(in_data_reg_69),
	.src_valid1(src_valid1),
	.out_byte_cnt_reg_2(out_byte_cnt_reg_2),
	.out_uncomp_byte_cnt_reg_4(out_uncomp_byte_cnt_reg_4),
	.out_uncomp_byte_cnt_reg_3(out_uncomp_byte_cnt_reg_3),
	.out_uncomp_byte_cnt_reg_2(out_uncomp_byte_cnt_reg_2),
	.out_uncomp_byte_cnt_reg_5(out_uncomp_byte_cnt_reg_5),
	.out_uncomp_byte_cnt_reg_6(out_uncomp_byte_cnt_reg_6),
	.sink0_endofpacket(src_payload_0),
	.in_data_reg_105(in_data_reg_105),
	.in_data_reg_106(in_data_reg_106),
	.in_data_reg_107(in_data_reg_107),
	.in_data_reg_108(in_data_reg_108),
	.in_data_reg_109(in_data_reg_109),
	.in_data_reg_110(in_data_reg_110),
	.in_data_reg_111(in_data_reg_111),
	.in_data_reg_112(in_data_reg_112),
	.in_data_reg_113(in_data_reg_113),
	.in_data_reg_114(in_data_reg_114),
	.in_data_reg_115(in_data_reg_115),
	.in_data_reg_116(in_data_reg_116),
	.Selector3(Selector3),
	.Selector10(Selector10),
	.base_address_3(base_address_3),
	.Selector4(Selector4),
	.Selector11(Selector11),
	.base_address_2(base_address_2),
	.Selector5(Selector5),
	.Selector12(Selector12),
	.out_data_1(out_data_1),
	.out_data_0(out_data_0),
	.Selector6(Selector6),
	.Selector13(Selector13),
	.clk_clk(clk_clk));

endmodule

module spw_babasu_altera_merlin_burst_adapter_13_1_14 (
	h2f_ARADDR_0,
	h2f_ARADDR_1,
	h2f_ARADDR_2,
	h2f_ARADDR_3,
	h2f_ARLEN_0,
	nxt_in_ready,
	in_ready_hold,
	stateST_COMP_TRANS,
	out_valid_reg1,
	in_narrow_reg1,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	in_data_reg_68,
	cp_ready,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready1,
	sink0_data,
	Equal15,
	altera_reset_synchronizer_int_chain_out,
	in_data_reg_0,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	in_data_reg_1,
	in_data_reg_2,
	in_data_reg_3,
	in_data_reg_4,
	in_data_reg_5,
	in_data_reg_6,
	Add2,
	Add21,
	Add22,
	Add23,
	write_cp_data_77,
	write_cp_data_78,
	write_cp_data_75,
	write_cp_data_74,
	write_cp_data_76,
	WideNor0,
	nxt_out_eop,
	Equal151,
	src15_valid,
	src_valid,
	cp_ready1,
	in_data_reg_69,
	src_valid1,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_6,
	sink0_endofpacket,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	Selector3,
	Selector10,
	base_address_3,
	Selector4,
	Selector11,
	base_address_2,
	Selector5,
	Selector12,
	out_data_1,
	out_data_0,
	Selector6,
	Selector13,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARADDR_0;
input 	h2f_ARADDR_1;
input 	h2f_ARADDR_2;
input 	h2f_ARADDR_3;
input 	h2f_ARLEN_0;
output 	nxt_in_ready;
input 	in_ready_hold;
output 	stateST_COMP_TRANS;
output 	out_valid_reg1;
output 	in_narrow_reg1;
output 	in_byteen_reg_3;
output 	in_byteen_reg_2;
output 	in_byteen_reg_1;
output 	in_byteen_reg_0;
output 	in_data_reg_68;
input 	cp_ready;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready1;
input 	[128:0] sink0_data;
input 	Equal15;
input 	altera_reset_synchronizer_int_chain_out;
output 	in_data_reg_0;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
output 	in_data_reg_1;
output 	in_data_reg_2;
output 	in_data_reg_3;
output 	in_data_reg_4;
output 	in_data_reg_5;
output 	in_data_reg_6;
input 	Add2;
input 	Add21;
input 	Add22;
input 	Add23;
input 	write_cp_data_77;
input 	write_cp_data_78;
input 	write_cp_data_75;
input 	write_cp_data_74;
input 	write_cp_data_76;
input 	WideNor0;
output 	nxt_out_eop;
input 	Equal151;
input 	src15_valid;
input 	src_valid;
input 	cp_ready1;
output 	in_data_reg_69;
input 	src_valid1;
output 	out_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_6;
input 	sink0_endofpacket;
output 	in_data_reg_105;
output 	in_data_reg_106;
output 	in_data_reg_107;
output 	in_data_reg_108;
output 	in_data_reg_109;
output 	in_data_reg_110;
output 	in_data_reg_111;
output 	in_data_reg_112;
output 	in_data_reg_113;
output 	in_data_reg_114;
output 	in_data_reg_115;
output 	in_data_reg_116;
input 	Selector3;
input 	Selector10;
input 	base_address_3;
input 	Selector4;
input 	Selector11;
input 	base_address_2;
input 	Selector5;
input 	Selector12;
input 	out_data_1;
input 	out_data_0;
input 	Selector6;
input 	Selector13;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \align_address_to_size|LessThan0~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt[4]~1_combout ;
wire \nxt_uncomp_subburst_byte_cnt[3]~2_combout ;
wire \Add4~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt[5]~3_combout ;
wire \nxt_uncomp_subburst_byte_cnt[2]~4_combout ;
wire \nxt_uncomp_subburst_byte_cnt[6]~5_combout ;
wire \WideOr0~combout ;
wire \in_valid~combout ;
wire \Selector0~0_combout ;
wire \load_next_out_cmd~combout ;
wire \state.ST_IDLE~q ;
wire \Selector2~0_combout ;
wire \Selector2~1_combout ;
wire \Selector2~2_combout ;
wire \state.ST_UNCOMP_TRANS~q ;
wire \Selector1~2_combout ;
wire \Selector1~0_combout ;
wire \Selector1~3_combout ;
wire \int_bytes_remaining_reg[5]~q ;
wire \d0_int_bytes_remaining[2]~4_combout ;
wire \d0_int_bytes_remaining[2]~5_combout ;
wire \int_bytes_remaining_reg[2]~q ;
wire \d0_int_bytes_remaining[3]~6_combout ;
wire \d0_int_bytes_remaining[3]~7_combout ;
wire \int_bytes_remaining_reg[3]~q ;
wire \Add1~1_combout ;
wire \d0_int_bytes_remaining[4]~8_combout ;
wire \int_bytes_remaining_reg[4]~q ;
wire \Add1~0_combout ;
wire \d0_int_bytes_remaining[5]~0_combout ;
wire \d0_int_bytes_remaining[5]~1_combout ;
wire \int_bytes_remaining_reg[6]~q ;
wire \d0_int_bytes_remaining[6]~2_combout ;
wire \d0_int_bytes_remaining[6]~3_combout ;
wire \Equal0~0_combout ;
wire \new_burst_reg~0_combout ;
wire \new_burst_reg~q ;
wire \Selector1~1_combout ;
wire \WideNor0~0_combout ;
wire \NON_PIPELINED_INPUTS.load_next_cmd~combout ;
wire \in_bytecount_reg_zero~q ;
wire \nxt_out_valid~0_combout ;
wire \LessThan0~0_combout ;
wire \Selector3~0_combout ;
wire \in_size_reg[0]~q ;
wire \in_size_reg[2]~q ;
wire \in_size_reg[1]~q ;
wire \ShiftLeft0~0_combout ;
wire \ShiftLeft0~1_combout ;
wire \int_byte_cnt_narrow_reg[3]~q ;
wire \ShiftLeft0~2_combout ;
wire \int_byte_cnt_narrow_reg[2]~q ;
wire \ShiftLeft0~3_combout ;
wire \ShiftLeft0~4_combout ;
wire \int_byte_cnt_narrow_reg[1]~q ;
wire \int_byte_cnt_narrow_reg[0]~q ;
wire \Add0~13_sumout ;
wire \d0_int_nxt_addr[0]~3_combout ;
wire \in_burstwrap_reg[0]~q ;
wire \nxt_addr[0]~0_combout ;
wire \int_nxt_addr_reg[0]~q ;
wire \d0_int_nxt_addr[0]~4_combout ;
wire \int_nxt_addr_reg_dly[0]~q ;
wire \Add0~14 ;
wire \Add0~9_sumout ;
wire \in_burstwrap_reg[1]~q ;
wire \nxt_addr[1]~4_combout ;
wire \int_nxt_addr_reg[1]~q ;
wire \d0_int_nxt_addr[1]~7_combout ;
wire \d0_int_nxt_addr[1]~2_combout ;
wire \int_nxt_addr_reg_dly[1]~q ;
wire \Add0~10 ;
wire \Add0~6 ;
wire \Add0~1_sumout ;
wire \in_burstwrap_reg[3]~q ;
wire \nxt_addr[3]~12_combout ;
wire \int_nxt_addr_reg[3]~q ;
wire \d0_int_nxt_addr[3]~5_combout ;
wire \d0_int_nxt_addr[3]~0_combout ;
wire \Add0~5_sumout ;
wire \in_burstwrap_reg[2]~q ;
wire \nxt_addr[2]~8_combout ;
wire \int_nxt_addr_reg[2]~q ;
wire \d0_int_nxt_addr[2]~6_combout ;
wire \d0_int_nxt_addr[2]~1_combout ;
wire \in_eop_reg~q ;


spw_babasu_altera_merlin_address_alignment_15 align_address_to_size(
	.new_burst_reg(\new_burst_reg~q ),
	.src_data_86(sink0_data[86]),
	.in_size_reg_0(\in_size_reg[0]~q ),
	.ShiftLeft0(\ShiftLeft0~3_combout ),
	.LessThan0(\align_address_to_size|LessThan0~0_combout ));

cyclonev_lcell_comb \nxt_in_ready~1 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!in_ready_hold),
	.datac(!out_valid_reg1),
	.datad(!cp_ready),
	.datae(!stateST_COMP_TRANS),
	.dataf(!\new_burst_reg~q ),
	.datag(!stateST_UNCOMP_WR_SUBBURST),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~1 .extended_lut = "on";
defparam \nxt_in_ready~1 .lut_mask = 64'h2020F0F02020F0FF;
defparam \nxt_in_ready~1 .shared_arith = "off";

dffeas \state.ST_COMP_TRANS (
	.clk(clk_clk),
	.d(\Selector1~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_COMP_TRANS),
	.prn(vcc));
defparam \state.ST_COMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_COMP_TRANS .power_up = "low";

dffeas out_valid_reg(
	.clk(clk_clk),
	.d(\nxt_out_valid~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_valid_reg1),
	.prn(vcc));
defparam out_valid_reg.is_wysiwyg = "true";
defparam out_valid_reg.power_up = "low";

dffeas in_narrow_reg(
	.clk(clk_clk),
	.d(\LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_narrow_reg1),
	.prn(vcc));
defparam in_narrow_reg.is_wysiwyg = "true";
defparam in_narrow_reg.power_up = "low";

dffeas \in_byteen_reg[3] (
	.clk(clk_clk),
	.d(sink0_data[35]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_3),
	.prn(vcc));
defparam \in_byteen_reg[3] .is_wysiwyg = "true";
defparam \in_byteen_reg[3] .power_up = "low";

dffeas \in_byteen_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[34]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_2),
	.prn(vcc));
defparam \in_byteen_reg[2] .is_wysiwyg = "true";
defparam \in_byteen_reg[2] .power_up = "low";

dffeas \in_byteen_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[33]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_1),
	.prn(vcc));
defparam \in_byteen_reg[1] .is_wysiwyg = "true";
defparam \in_byteen_reg[1] .power_up = "low";

dffeas \in_byteen_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[32]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_0),
	.prn(vcc));
defparam \in_byteen_reg[0] .is_wysiwyg = "true";
defparam \in_byteen_reg[0] .power_up = "low";

dffeas \in_data_reg[68] (
	.clk(clk_clk),
	.d(sink0_data[68]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_68),
	.prn(vcc));
defparam \in_data_reg[68] .is_wysiwyg = "true";
defparam \in_data_reg[68] .power_up = "low";

dffeas \state.ST_UNCOMP_WR_SUBBURST (
	.clk(clk_clk),
	.d(\Selector3~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_UNCOMP_WR_SUBBURST),
	.prn(vcc));
defparam \state.ST_UNCOMP_WR_SUBBURST .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_WR_SUBBURST .power_up = "low";

cyclonev_lcell_comb \nxt_in_ready~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!out_valid_reg1),
	.datac(!cp_ready),
	.datad(!\state.ST_UNCOMP_TRANS~q ),
	.datae(!stateST_UNCOMP_WR_SUBBURST),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~0 .extended_lut = "off";
defparam \nxt_in_ready~0 .lut_mask = 64'h008A8A8A008A8A8A;
defparam \nxt_in_ready~0 .shared_arith = "off";

dffeas \in_data_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[0]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_0),
	.prn(vcc));
defparam \in_data_reg[0] .is_wysiwyg = "true";
defparam \in_data_reg[0] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[3] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[3]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_3),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[3] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[2] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[2]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_2),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[2] .power_up = "low";

dffeas \in_data_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[1]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_1),
	.prn(vcc));
defparam \in_data_reg[1] .is_wysiwyg = "true";
defparam \in_data_reg[1] .power_up = "low";

dffeas \in_data_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[2]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_2),
	.prn(vcc));
defparam \in_data_reg[2] .is_wysiwyg = "true";
defparam \in_data_reg[2] .power_up = "low";

dffeas \in_data_reg[3] (
	.clk(clk_clk),
	.d(sink0_data[3]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_3),
	.prn(vcc));
defparam \in_data_reg[3] .is_wysiwyg = "true";
defparam \in_data_reg[3] .power_up = "low";

dffeas \in_data_reg[4] (
	.clk(clk_clk),
	.d(sink0_data[4]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_4),
	.prn(vcc));
defparam \in_data_reg[4] .is_wysiwyg = "true";
defparam \in_data_reg[4] .power_up = "low";

dffeas \in_data_reg[5] (
	.clk(clk_clk),
	.d(sink0_data[5]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_5),
	.prn(vcc));
defparam \in_data_reg[5] .is_wysiwyg = "true";
defparam \in_data_reg[5] .power_up = "low";

dffeas \in_data_reg[6] (
	.clk(clk_clk),
	.d(sink0_data[6]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_6),
	.prn(vcc));
defparam \in_data_reg[6] .is_wysiwyg = "true";
defparam \in_data_reg[6] .power_up = "low";

cyclonev_lcell_comb \nxt_out_eop~0 (
	.dataa(!\in_eop_reg~q ),
	.datab(!stateST_COMP_TRANS),
	.datac(!\new_burst_reg~q ),
	.datad(!cp_ready),
	.datae(!\in_bytecount_reg_zero~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_out_eop),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_eop~0 .extended_lut = "off";
defparam \nxt_out_eop~0 .lut_mask = 64'h4447774744477747;
defparam \nxt_out_eop~0 .shared_arith = "off";

dffeas \in_data_reg[69] (
	.clk(clk_clk),
	.d(sink0_data[69]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_69),
	.prn(vcc));
defparam \in_data_reg[69] .is_wysiwyg = "true";
defparam \in_data_reg[69] .power_up = "low";

dffeas \out_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[4] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[4]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_4),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[4] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[4] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[3] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[3]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_3),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[3] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[3] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[2]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[5] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[5]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_5),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[5] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[5] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[6] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[6]~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_6),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[6] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[6] .power_up = "low";

dffeas \in_data_reg[105] (
	.clk(clk_clk),
	.d(sink0_data[105]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_105),
	.prn(vcc));
defparam \in_data_reg[105] .is_wysiwyg = "true";
defparam \in_data_reg[105] .power_up = "low";

dffeas \in_data_reg[106] (
	.clk(clk_clk),
	.d(sink0_data[106]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_106),
	.prn(vcc));
defparam \in_data_reg[106] .is_wysiwyg = "true";
defparam \in_data_reg[106] .power_up = "low";

dffeas \in_data_reg[107] (
	.clk(clk_clk),
	.d(sink0_data[107]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_107),
	.prn(vcc));
defparam \in_data_reg[107] .is_wysiwyg = "true";
defparam \in_data_reg[107] .power_up = "low";

dffeas \in_data_reg[108] (
	.clk(clk_clk),
	.d(sink0_data[108]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_108),
	.prn(vcc));
defparam \in_data_reg[108] .is_wysiwyg = "true";
defparam \in_data_reg[108] .power_up = "low";

dffeas \in_data_reg[109] (
	.clk(clk_clk),
	.d(sink0_data[109]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_109),
	.prn(vcc));
defparam \in_data_reg[109] .is_wysiwyg = "true";
defparam \in_data_reg[109] .power_up = "low";

dffeas \in_data_reg[110] (
	.clk(clk_clk),
	.d(sink0_data[110]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_110),
	.prn(vcc));
defparam \in_data_reg[110] .is_wysiwyg = "true";
defparam \in_data_reg[110] .power_up = "low";

dffeas \in_data_reg[111] (
	.clk(clk_clk),
	.d(sink0_data[111]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_111),
	.prn(vcc));
defparam \in_data_reg[111] .is_wysiwyg = "true";
defparam \in_data_reg[111] .power_up = "low";

dffeas \in_data_reg[112] (
	.clk(clk_clk),
	.d(sink0_data[112]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_112),
	.prn(vcc));
defparam \in_data_reg[112] .is_wysiwyg = "true";
defparam \in_data_reg[112] .power_up = "low";

dffeas \in_data_reg[113] (
	.clk(clk_clk),
	.d(sink0_data[113]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_113),
	.prn(vcc));
defparam \in_data_reg[113] .is_wysiwyg = "true";
defparam \in_data_reg[113] .power_up = "low";

dffeas \in_data_reg[114] (
	.clk(clk_clk),
	.d(sink0_data[114]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_114),
	.prn(vcc));
defparam \in_data_reg[114] .is_wysiwyg = "true";
defparam \in_data_reg[114] .power_up = "low";

dffeas \in_data_reg[115] (
	.clk(clk_clk),
	.d(sink0_data[115]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_115),
	.prn(vcc));
defparam \in_data_reg[115] .is_wysiwyg = "true";
defparam \in_data_reg[115] .power_up = "low";

dffeas \in_data_reg[116] (
	.clk(clk_clk),
	.d(sink0_data[116]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_116),
	.prn(vcc));
defparam \in_data_reg[116] .is_wysiwyg = "true";
defparam \in_data_reg[116] .power_up = "low";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt~0 (
	.dataa(!out_valid_reg1),
	.datab(!cp_ready),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt~0 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt~0 .lut_mask = 64'h1111111111111111;
defparam \nxt_uncomp_subburst_byte_cnt~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[4]~1 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!out_uncomp_byte_cnt_reg_3),
	.datae(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.dataf(!out_uncomp_byte_cnt_reg_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[4]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[4]~1 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[4]~1 .lut_mask = 64'h0F0FE44E0F0F4E4E;
defparam \nxt_uncomp_subburst_byte_cnt[4]~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[3]~2 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!out_uncomp_byte_cnt_reg_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[3]~2 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[3]~2 .lut_mask = 64'h0FE40F4E0FE40F4E;
defparam \nxt_uncomp_subburst_byte_cnt[3]~2 .shared_arith = "off";

cyclonev_lcell_comb \Add4~0 (
	.dataa(!out_uncomp_byte_cnt_reg_4),
	.datab(!out_uncomp_byte_cnt_reg_3),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add4~0 .extended_lut = "off";
defparam \Add4~0 .lut_mask = 64'h0800080008000800;
defparam \Add4~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[5]~3 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_5),
	.datae(!\Add4~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[5]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[5]~3 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[5]~3 .lut_mask = 64'h04FEAE5404FEAE54;
defparam \nxt_uncomp_subburst_byte_cnt[5]~3 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[2]~4 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[2]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[2]~4 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[2]~4 .lut_mask = 64'h0EF40EF40EF40EF4;
defparam \nxt_uncomp_subburst_byte_cnt[2]~4 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[6]~5 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_5),
	.datae(!\Add4~0_combout ),
	.dataf(!out_uncomp_byte_cnt_reg_6),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[6]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[6]~5 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[6]~5 .lut_mask = 64'h0404AE04FEFE54FE;
defparam \nxt_uncomp_subburst_byte_cnt[6]~5 .shared_arith = "off";

cyclonev_lcell_comb WideOr0(
	.dataa(!\nxt_uncomp_subburst_byte_cnt[4]~1_combout ),
	.datab(!\nxt_uncomp_subburst_byte_cnt[3]~2_combout ),
	.datac(!\nxt_uncomp_subburst_byte_cnt[5]~3_combout ),
	.datad(!\nxt_uncomp_subburst_byte_cnt[2]~4_combout ),
	.datae(!\nxt_uncomp_subburst_byte_cnt[6]~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr0.extended_lut = "off";
defparam WideOr0.lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam WideOr0.shared_arith = "off";

cyclonev_lcell_comb in_valid(
	.dataa(!in_ready_hold),
	.datab(!Equal15),
	.datac(!Equal151),
	.datad(!sink0_data[68]),
	.datae(!src15_valid),
	.dataf(!src_valid),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\in_valid~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam in_valid.extended_lut = "off";
defparam in_valid.lut_mask = 64'h0000000155555555;
defparam in_valid.shared_arith = "off";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!sink0_data[69]),
	.datab(!nxt_out_eop),
	.datac(!sink0_data[68]),
	.datad(!\in_valid~combout ),
	.datae(!\state.ST_IDLE~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'h005FCCFF005FCCFF;
defparam \Selector0~0 .shared_arith = "off";

cyclonev_lcell_comb load_next_out_cmd(
	.dataa(!out_valid_reg1),
	.datab(!cp_ready),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\load_next_out_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam load_next_out_cmd.extended_lut = "off";
defparam load_next_out_cmd.lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam load_next_out_cmd.shared_arith = "off";

dffeas \state.ST_IDLE (
	.clk(clk_clk),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_IDLE~q ),
	.prn(vcc));
defparam \state.ST_IDLE .is_wysiwyg = "true";
defparam \state.ST_IDLE .power_up = "low";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!nxt_out_eop),
	.datac(!stateST_UNCOMP_WR_SUBBURST),
	.datad(!\state.ST_IDLE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'h00EC00EC00EC00EC;
defparam \Selector2~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~1 (
	.dataa(!in_ready_hold),
	.datab(!Equal15),
	.datac(!Equal151),
	.datad(!sink0_data[68]),
	.datae(!src15_valid),
	.dataf(!\Selector2~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~1 .extended_lut = "off";
defparam \Selector2~1 .lut_mask = 64'h0000000100000000;
defparam \Selector2~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~2 (
	.dataa(!\WideOr0~combout ),
	.datab(!\Selector2~1_combout ),
	.datac(!\in_valid~combout ),
	.datad(!nxt_out_eop),
	.datae(!\state.ST_UNCOMP_TRANS~q ),
	.dataf(!sink0_data[69]),
	.datag(!stateST_UNCOMP_WR_SUBBURST),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~2 .extended_lut = "on";
defparam \Selector2~2 .lut_mask = 64'h3B33BB3F0A00AA00;
defparam \Selector2~2 .shared_arith = "off";

dffeas \state.ST_UNCOMP_TRANS (
	.clk(clk_clk),
	.d(\Selector2~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_UNCOMP_TRANS~q ),
	.prn(vcc));
defparam \state.ST_UNCOMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_TRANS .power_up = "low";

cyclonev_lcell_comb \Selector1~2 (
	.dataa(!in_ready_hold),
	.datab(!stateST_COMP_TRANS),
	.datac(!nxt_out_eop),
	.datad(!sink0_data[68]),
	.datae(gnd),
	.dataf(!src_valid),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~2 .extended_lut = "off";
defparam \Selector1~2 .lut_mask = 64'h3030303031303130;
defparam \Selector1~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!nxt_out_eop),
	.datac(!\state.ST_UNCOMP_TRANS~q ),
	.datad(!stateST_UNCOMP_WR_SUBBURST),
	.datae(!\state.ST_IDLE~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'h0000A8880000A888;
defparam \Selector1~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~3 (
	.dataa(!in_ready_hold),
	.datab(!sink0_data[69]),
	.datac(!src_valid),
	.datad(!src_valid1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~3 .extended_lut = "off";
defparam \Selector1~3 .lut_mask = 64'h0111011101110111;
defparam \Selector1~3 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[5] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[5]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[5]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[5] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[5] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[2]~4 (
	.dataa(!h2f_ARLEN_0),
	.datab(!sink0_data[69]),
	.datac(!sink0_data[68]),
	.datad(!write_cp_data_74),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[2]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[2]~4 .extended_lut = "off";
defparam \d0_int_bytes_remaining[2]~4 .lut_mask = 64'h2F222F222F222F22;
defparam \d0_int_bytes_remaining[2]~4 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[2]~5 (
	.dataa(!\new_burst_reg~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\int_bytes_remaining_reg[2]~q ),
	.datad(!\d0_int_bytes_remaining[2]~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[2]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[2]~5 .extended_lut = "off";
defparam \d0_int_bytes_remaining[2]~5 .lut_mask = 64'h287D287D287D287D;
defparam \d0_int_bytes_remaining[2]~5 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[2] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[2]~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[2]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[2] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[3]~6 (
	.dataa(!sink0_data[69]),
	.datab(!sink0_data[68]),
	.datac(!write_cp_data_75),
	.datad(!Add2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[3]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[3]~6 .extended_lut = "off";
defparam \d0_int_bytes_remaining[3]~6 .lut_mask = 64'h0357035703570357;
defparam \d0_int_bytes_remaining[3]~6 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[3]~7 (
	.dataa(!\new_burst_reg~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\int_bytes_remaining_reg[2]~q ),
	.datad(!\int_bytes_remaining_reg[3]~q ),
	.datae(!\d0_int_bytes_remaining[3]~6_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[3]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[3]~7 .extended_lut = "off";
defparam \d0_int_bytes_remaining[3]~7 .lut_mask = 64'h208A75DF208A75DF;
defparam \d0_int_bytes_remaining[3]~7 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[3] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[3]~7_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[3]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[3] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[3] .power_up = "low";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!out_byte_cnt_reg_2),
	.datab(!\int_bytes_remaining_reg[2]~q ),
	.datac(!\int_bytes_remaining_reg[3]~q ),
	.datad(!\int_bytes_remaining_reg[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'hBF40BF40BF40BF40;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[4]~8 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!sink0_data[68]),
	.datad(!write_cp_data_76),
	.datae(!Add21),
	.dataf(!\Add1~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[4]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[4]~8 .extended_lut = "off";
defparam \d0_int_bytes_remaining[4]~8 .lut_mask = 64'hCCCFDDDF00031113;
defparam \d0_int_bytes_remaining[4]~8 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[4] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[4]~8_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[4]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[4] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[4] .power_up = "low";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!out_byte_cnt_reg_2),
	.datab(!\int_bytes_remaining_reg[2]~q ),
	.datac(!\int_bytes_remaining_reg[3]~q ),
	.datad(!\int_bytes_remaining_reg[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h4000400040004000;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[5]~0 (
	.dataa(!sink0_data[69]),
	.datab(!sink0_data[68]),
	.datac(!write_cp_data_77),
	.datad(!Add22),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[5]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[5]~0 .extended_lut = "off";
defparam \d0_int_bytes_remaining[5]~0 .lut_mask = 64'h0357035703570357;
defparam \d0_int_bytes_remaining[5]~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[5]~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\int_bytes_remaining_reg[5]~q ),
	.datac(!\Add1~0_combout ),
	.datad(!\d0_int_bytes_remaining[5]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[5]~1 .extended_lut = "off";
defparam \d0_int_bytes_remaining[5]~1 .lut_mask = 64'h287D287D287D287D;
defparam \d0_int_bytes_remaining[5]~1 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[6] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[6]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[6]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[6] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[6] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[6]~2 (
	.dataa(!sink0_data[69]),
	.datab(!sink0_data[68]),
	.datac(!write_cp_data_78),
	.datad(!Add23),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[6]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[6]~2 .extended_lut = "off";
defparam \d0_int_bytes_remaining[6]~2 .lut_mask = 64'h0357035703570357;
defparam \d0_int_bytes_remaining[6]~2 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[6]~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\int_bytes_remaining_reg[5]~q ),
	.datac(!\Add1~0_combout ),
	.datad(!\int_bytes_remaining_reg[6]~q ),
	.datae(!\d0_int_bytes_remaining[6]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[6]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[6]~3 .extended_lut = "off";
defparam \d0_int_bytes_remaining[6]~3 .lut_mask = 64'h08A25DF708A25DF7;
defparam \d0_int_bytes_remaining[6]~3 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!\d0_int_bytes_remaining[2]~5_combout ),
	.datab(!\d0_int_bytes_remaining[3]~7_combout ),
	.datac(!\d0_int_bytes_remaining[4]~8_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'h4040404040404040;
defparam \Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \new_burst_reg~0 (
	.dataa(!\Selector1~2_combout ),
	.datab(!\Selector1~0_combout ),
	.datac(!\Selector1~3_combout ),
	.datad(!\d0_int_bytes_remaining[5]~1_combout ),
	.datae(!\d0_int_bytes_remaining[6]~3_combout ),
	.dataf(!\Equal0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\new_burst_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \new_burst_reg~0 .extended_lut = "off";
defparam \new_burst_reg~0 .lut_mask = 64'hA2A2A2A2FFA2A2A2;
defparam \new_burst_reg~0 .shared_arith = "off";

dffeas new_burst_reg(
	.clk(clk_clk),
	.d(\new_burst_reg~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\new_burst_reg~q ),
	.prn(vcc));
defparam new_burst_reg.is_wysiwyg = "true";
defparam new_burst_reg.power_up = "low";

cyclonev_lcell_comb \Selector1~1 (
	.dataa(!sink0_data[69]),
	.datab(!stateST_COMP_TRANS),
	.datac(!nxt_out_eop),
	.datad(!sink0_data[68]),
	.datae(!\in_valid~combout ),
	.dataf(!\Selector1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~1 .extended_lut = "off";
defparam \Selector1~1 .lut_mask = 64'h3030777530303330;
defparam \Selector1~1 .shared_arith = "off";

cyclonev_lcell_comb \WideNor0~0 (
	.dataa(!sink0_data[69]),
	.datab(!sink0_data[68]),
	.datac(!WideNor0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideNor0~0 .extended_lut = "off";
defparam \WideNor0~0 .lut_mask = 64'h8A8A8A8A8A8A8A8A;
defparam \WideNor0~0 .shared_arith = "off";

cyclonev_lcell_comb \NON_PIPELINED_INPUTS.load_next_cmd (
	.dataa(!in_ready_hold),
	.datab(!nxt_in_ready1),
	.datac(!nxt_in_ready),
	.datad(!src_valid),
	.datae(!src_valid1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \NON_PIPELINED_INPUTS.load_next_cmd .extended_lut = "off";
defparam \NON_PIPELINED_INPUTS.load_next_cmd .lut_mask = 64'h0015151500151515;
defparam \NON_PIPELINED_INPUTS.load_next_cmd .shared_arith = "off";

dffeas in_bytecount_reg_zero(
	.clk(clk_clk),
	.d(\WideNor0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_bytecount_reg_zero~q ),
	.prn(vcc));
defparam in_bytecount_reg_zero.is_wysiwyg = "true";
defparam in_bytecount_reg_zero.power_up = "low";

cyclonev_lcell_comb \nxt_out_valid~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!\new_burst_reg~q ),
	.datac(!\in_bytecount_reg_zero~q ),
	.datad(!\in_valid~combout ),
	.datae(!cp_ready1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_valid~0 .extended_lut = "off";
defparam \nxt_out_valid~0 .lut_mask = 64'h50FF44FF50FF44FF;
defparam \nxt_out_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!sink0_data[87]),
	.datab(!sink0_data[88]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h8888888888888888;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~0 (
	.dataa(!nxt_out_eop),
	.datab(!\state.ST_UNCOMP_TRANS~q ),
	.datac(!stateST_UNCOMP_WR_SUBBURST),
	.datad(!\WideOr0~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'h002A002A002A002A;
defparam \Selector3~0 .shared_arith = "off";

dffeas \in_size_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[86]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[0]~q ),
	.prn(vcc));
defparam \in_size_reg[0] .is_wysiwyg = "true";
defparam \in_size_reg[0] .power_up = "low";

dffeas \in_size_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[88]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[2]~q ),
	.prn(vcc));
defparam \in_size_reg[2] .is_wysiwyg = "true";
defparam \in_size_reg[2] .power_up = "low";

dffeas \in_size_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[87]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[1]~q ),
	.prn(vcc));
defparam \in_size_reg[1] .is_wysiwyg = "true";
defparam \in_size_reg[1] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[87]),
	.datac(!sink0_data[88]),
	.datad(!\in_size_reg[2]~q ),
	.datae(!\in_size_reg[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~0 .extended_lut = "off";
defparam \ShiftLeft0~0 .lut_mask = 64'h1010BA101010BA10;
defparam \ShiftLeft0~0 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~1 .extended_lut = "off";
defparam \ShiftLeft0~1 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~1 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[3] (
	.clk(clk_clk),
	.d(\ShiftLeft0~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[3]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[3] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[3] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~2 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~2 .extended_lut = "off";
defparam \ShiftLeft0~2 .lut_mask = 64'h00E400E400E400E4;
defparam \ShiftLeft0~2 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[2] (
	.clk(clk_clk),
	.d(\ShiftLeft0~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[2]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[2] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[2] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[87]),
	.datac(!sink0_data[88]),
	.datad(!\in_size_reg[2]~q ),
	.datae(!\in_size_reg[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~3 .extended_lut = "off";
defparam \ShiftLeft0~3 .lut_mask = 64'hEA404040EA404040;
defparam \ShiftLeft0~3 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~4 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~4 .extended_lut = "off";
defparam \ShiftLeft0~4 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~4 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[1] (
	.clk(clk_clk),
	.d(\ShiftLeft0~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[1]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[1] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[1] .power_up = "low";

dffeas \int_byte_cnt_narrow_reg[0] (
	.clk(clk_clk),
	.d(\align_address_to_size|LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[0]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[0] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[0] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[0]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~3 (
	.dataa(!h2f_ARADDR_0),
	.datab(!sink0_data[69]),
	.datac(!sink0_data[68]),
	.datad(!out_data_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~3 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~3 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[0]~3 .shared_arith = "off";

dffeas \in_burstwrap_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[79]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[0]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[0] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[0] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[0]~0 (
	.dataa(!Selector13),
	.datab(!Selector6),
	.datac(!sink0_data[68]),
	.datad(!sink0_data[69]),
	.datae(!\new_burst_reg~q ),
	.dataf(!\d0_int_nxt_addr[0]~4_combout ),
	.datag(!\in_burstwrap_reg[0]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[0]~0 .extended_lut = "on";
defparam \nxt_addr[0]~0 .lut_mask = 64'h00000000F0F0FCA8;
defparam \nxt_addr[0]~0 .shared_arith = "off";

dffeas \int_nxt_addr_reg[0] (
	.clk(clk_clk),
	.d(\nxt_addr[0]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[0] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~4 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\Add0~13_sumout ),
	.datac(!\align_address_to_size|LessThan0~0_combout ),
	.datad(!\d0_int_nxt_addr[0]~3_combout ),
	.datae(!\int_nxt_addr_reg[0]~q ),
	.dataf(!\in_burstwrap_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~4 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~4 .lut_mask = 64'h0005AAAF2227AAAF;
defparam \d0_int_nxt_addr[0]~4 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[0] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[0]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[0] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[1]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[1]~q ),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \in_burstwrap_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[80]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[1]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[1] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[1] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[1]~4 (
	.dataa(!Selector12),
	.datab(!Selector5),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!\new_burst_reg~q ),
	.dataf(!\d0_int_nxt_addr[1]~2_combout ),
	.datag(!\in_burstwrap_reg[1]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[1]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[1]~4 .extended_lut = "on";
defparam \nxt_addr[1]~4 .lut_mask = 64'h00000000F0F0FAC8;
defparam \nxt_addr[1]~4 .shared_arith = "off";

dffeas \int_nxt_addr_reg[1] (
	.clk(clk_clk),
	.d(\nxt_addr[1]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[1] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~7 (
	.dataa(!h2f_ARADDR_1),
	.datab(!sink0_data[69]),
	.datac(!sink0_data[68]),
	.datad(!out_data_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~7 .extended_lut = "off";
defparam \d0_int_nxt_addr[1]~7 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[1]~7 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~2 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\Add0~9_sumout ),
	.datac(!\in_burstwrap_reg[1]~q ),
	.datad(!\int_nxt_addr_reg[1]~q ),
	.datae(!\ShiftLeft0~3_combout ),
	.dataf(!\d0_int_nxt_addr[1]~7_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~2 .extended_lut = "off";
defparam \d0_int_nxt_addr[1]~2 .lut_mask = 64'h02AA02AA02AA57FF;
defparam \d0_int_nxt_addr[1]~2 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[1] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[1]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[1] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_2),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[2]~q ),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[3]~q ),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

dffeas \in_burstwrap_reg[3] (
	.clk(clk_clk),
	.d(sink0_data[82]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[3]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[3] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[3] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[3]~12 (
	.dataa(!Selector10),
	.datab(!Selector3),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!\new_burst_reg~q ),
	.dataf(!\d0_int_nxt_addr[3]~0_combout ),
	.datag(!\in_burstwrap_reg[3]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[3]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[3]~12 .extended_lut = "on";
defparam \nxt_addr[3]~12 .lut_mask = 64'h00000000F0F0FAC8;
defparam \nxt_addr[3]~12 .shared_arith = "off";

dffeas \int_nxt_addr_reg[3] (
	.clk(clk_clk),
	.d(\nxt_addr[3]~12_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[3]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[3] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~5 (
	.dataa(!\Add0~1_sumout ),
	.datab(!\in_burstwrap_reg[3]~q ),
	.datac(!\int_nxt_addr_reg[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~5 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~5 .lut_mask = 64'hE0E0E0E0E0E0E0E0;
defparam \d0_int_nxt_addr[3]~5 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!h2f_ARADDR_3),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!base_address_3),
	.dataf(!\d0_int_nxt_addr[3]~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~0 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~0 .lut_mask = 64'hABABABFF01010155;
defparam \d0_int_nxt_addr[3]~0 .shared_arith = "off";

dffeas \in_burstwrap_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[81]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[2]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[2] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[2] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[2]~8 (
	.dataa(!Selector11),
	.datab(!Selector4),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!\new_burst_reg~q ),
	.dataf(!\d0_int_nxt_addr[2]~1_combout ),
	.datag(!\in_burstwrap_reg[2]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[2]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[2]~8 .extended_lut = "on";
defparam \nxt_addr[2]~8 .lut_mask = 64'h00000000F0F0FAC8;
defparam \nxt_addr[2]~8 .shared_arith = "off";

dffeas \int_nxt_addr_reg[2] (
	.clk(clk_clk),
	.d(\nxt_addr[2]~8_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[2]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~6 (
	.dataa(!\Add0~5_sumout ),
	.datab(!\in_burstwrap_reg[2]~q ),
	.datac(!\int_nxt_addr_reg[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~6 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~6 .lut_mask = 64'hE0E0E0E0E0E0E0E0;
defparam \d0_int_nxt_addr[2]~6 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!h2f_ARADDR_2),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!base_address_2),
	.dataf(!\d0_int_nxt_addr[2]~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~1 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~1 .lut_mask = 64'hABABABFF01010155;
defparam \d0_int_nxt_addr[2]~1 .shared_arith = "off";

dffeas in_eop_reg(
	.clk(clk_clk),
	.d(sink0_endofpacket),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_eop_reg~q ),
	.prn(vcc));
defparam in_eop_reg.is_wysiwyg = "true";
defparam in_eop_reg.power_up = "low";

endmodule

module spw_babasu_altera_merlin_address_alignment_15 (
	new_burst_reg,
	src_data_86,
	in_size_reg_0,
	ShiftLeft0,
	LessThan0)/* synthesis synthesis_greybox=0 */;
input 	new_burst_reg;
input 	src_data_86;
input 	in_size_reg_0;
input 	ShiftLeft0;
output 	LessThan0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!new_burst_reg),
	.datab(!src_data_86),
	.datac(!in_size_reg_0),
	.datad(!ShiftLeft0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan0),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h00E400E400E400E4;
defparam \LessThan0~0 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_burst_adapter_15 (
	h2f_ARADDR_0,
	h2f_ARADDR_1,
	h2f_ARADDR_2,
	h2f_ARADDR_3,
	h2f_ARBURST_0,
	h2f_ARBURST_1,
	h2f_ARID_0,
	h2f_ARID_1,
	h2f_ARID_2,
	h2f_ARID_3,
	h2f_ARID_4,
	h2f_ARID_5,
	h2f_ARID_6,
	h2f_ARID_7,
	h2f_ARID_8,
	h2f_ARID_9,
	h2f_ARID_10,
	h2f_ARID_11,
	h2f_ARLEN_0,
	Add5,
	Add51,
	in_ready_hold,
	in_data_reg_69,
	stateST_COMP_TRANS,
	mem_used_1,
	in_narrow_reg,
	cp_ready,
	nxt_in_ready,
	out_valid_reg,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready1,
	saved_grant_1,
	altera_reset_synchronizer_int_chain_out,
	Decoder1,
	Add2,
	Add21,
	Add22,
	Add23,
	nxt_in_ready2,
	src_valid,
	nxt_out_eop,
	out_byte_cnt_reg_2,
	cp_ready1,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_6,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	Selector10,
	Selector101,
	Selector11,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	Selector12,
	src_payload,
	src_payload1,
	src_payload2,
	Selector13,
	nxt_out_burstwrap_1,
	nxt_addr_2,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARADDR_0;
input 	h2f_ARADDR_1;
input 	h2f_ARADDR_2;
input 	h2f_ARADDR_3;
input 	h2f_ARBURST_0;
input 	h2f_ARBURST_1;
input 	h2f_ARID_0;
input 	h2f_ARID_1;
input 	h2f_ARID_2;
input 	h2f_ARID_3;
input 	h2f_ARID_4;
input 	h2f_ARID_5;
input 	h2f_ARID_6;
input 	h2f_ARID_7;
input 	h2f_ARID_8;
input 	h2f_ARID_9;
input 	h2f_ARID_10;
input 	h2f_ARID_11;
input 	h2f_ARLEN_0;
input 	Add5;
input 	Add51;
input 	in_ready_hold;
output 	in_data_reg_69;
output 	stateST_COMP_TRANS;
input 	mem_used_1;
output 	in_narrow_reg;
input 	cp_ready;
output 	nxt_in_ready;
output 	out_valid_reg;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready1;
input 	saved_grant_1;
input 	altera_reset_synchronizer_int_chain_out;
input 	Decoder1;
input 	Add2;
input 	Add21;
input 	Add22;
input 	Add23;
output 	nxt_in_ready2;
input 	src_valid;
output 	nxt_out_eop;
output 	out_byte_cnt_reg_2;
input 	cp_ready1;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_6;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_4;
output 	in_data_reg_105;
output 	in_data_reg_106;
output 	in_data_reg_107;
output 	in_data_reg_108;
output 	in_data_reg_109;
output 	in_data_reg_110;
output 	in_data_reg_111;
output 	in_data_reg_112;
output 	in_data_reg_113;
output 	in_data_reg_114;
output 	in_data_reg_115;
output 	in_data_reg_116;
input 	Selector10;
input 	Selector101;
input 	Selector11;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
input 	Selector12;
input 	src_payload;
input 	src_payload1;
input 	src_payload2;
input 	Selector13;
input 	nxt_out_burstwrap_1;
input 	nxt_addr_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



spw_babasu_altera_merlin_burst_adapter_13_1_15 \altera_merlin_burst_adapter_13_1.burst_adapter (
	.h2f_ARADDR_0(h2f_ARADDR_0),
	.h2f_ARADDR_1(h2f_ARADDR_1),
	.h2f_ARADDR_2(h2f_ARADDR_2),
	.h2f_ARADDR_3(h2f_ARADDR_3),
	.h2f_ARBURST_0(h2f_ARBURST_0),
	.h2f_ARBURST_1(h2f_ARBURST_1),
	.sink0_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,h2f_ARID_11,h2f_ARID_10,h2f_ARID_9,h2f_ARID_8,h2f_ARID_7,h2f_ARID_6,h2f_ARID_5,h2f_ARID_4,h2f_ARID_3,h2f_ARID_2,h2f_ARID_1,h2f_ARID_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_payload2,src_payload1,src_payload,gnd,gnd,gnd,
Selector101,Selector11,Selector12,Selector13,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,saved_grant_1,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.h2f_ARLEN_0(h2f_ARLEN_0),
	.Add5(Add5),
	.Add51(Add51),
	.in_ready_hold(in_ready_hold),
	.in_data_reg_69(in_data_reg_69),
	.stateST_COMP_TRANS(stateST_COMP_TRANS),
	.mem_used_1(mem_used_1),
	.in_narrow_reg1(in_narrow_reg),
	.cp_ready(cp_ready),
	.nxt_in_ready(nxt_in_ready),
	.out_valid_reg1(out_valid_reg),
	.stateST_UNCOMP_WR_SUBBURST(stateST_UNCOMP_WR_SUBBURST),
	.nxt_in_ready1(nxt_in_ready1),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.Decoder1(Decoder1),
	.Add2(Add2),
	.Add21(Add21),
	.Add22(Add22),
	.Add23(Add23),
	.nxt_in_ready2(nxt_in_ready2),
	.src_valid(src_valid),
	.nxt_out_eop(nxt_out_eop),
	.out_byte_cnt_reg_2(out_byte_cnt_reg_2),
	.cp_ready1(cp_ready1),
	.out_uncomp_byte_cnt_reg_3(out_uncomp_byte_cnt_reg_3),
	.out_uncomp_byte_cnt_reg_2(out_uncomp_byte_cnt_reg_2),
	.out_uncomp_byte_cnt_reg_6(out_uncomp_byte_cnt_reg_6),
	.out_uncomp_byte_cnt_reg_5(out_uncomp_byte_cnt_reg_5),
	.out_uncomp_byte_cnt_reg_4(out_uncomp_byte_cnt_reg_4),
	.in_data_reg_105(in_data_reg_105),
	.in_data_reg_106(in_data_reg_106),
	.in_data_reg_107(in_data_reg_107),
	.in_data_reg_108(in_data_reg_108),
	.in_data_reg_109(in_data_reg_109),
	.in_data_reg_110(in_data_reg_110),
	.in_data_reg_111(in_data_reg_111),
	.in_data_reg_112(in_data_reg_112),
	.in_data_reg_113(in_data_reg_113),
	.in_data_reg_114(in_data_reg_114),
	.in_data_reg_115(in_data_reg_115),
	.in_data_reg_116(in_data_reg_116),
	.Selector10(Selector10),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_3),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_2),
	.nxt_out_burstwrap_1(nxt_out_burstwrap_1),
	.nxt_addr_2(nxt_addr_2),
	.clk_clk(clk_clk));

endmodule

module spw_babasu_altera_merlin_burst_adapter_13_1_15 (
	h2f_ARADDR_0,
	h2f_ARADDR_1,
	h2f_ARADDR_2,
	h2f_ARADDR_3,
	h2f_ARBURST_0,
	h2f_ARBURST_1,
	sink0_data,
	h2f_ARLEN_0,
	Add5,
	Add51,
	in_ready_hold,
	in_data_reg_69,
	stateST_COMP_TRANS,
	mem_used_1,
	in_narrow_reg1,
	cp_ready,
	nxt_in_ready,
	out_valid_reg1,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready1,
	altera_reset_synchronizer_int_chain_out,
	Decoder1,
	Add2,
	Add21,
	Add22,
	Add23,
	nxt_in_ready2,
	src_valid,
	nxt_out_eop,
	out_byte_cnt_reg_2,
	cp_ready1,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_6,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	Selector10,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	nxt_out_burstwrap_1,
	nxt_addr_2,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARADDR_0;
input 	h2f_ARADDR_1;
input 	h2f_ARADDR_2;
input 	h2f_ARADDR_3;
input 	h2f_ARBURST_0;
input 	h2f_ARBURST_1;
input 	[128:0] sink0_data;
input 	h2f_ARLEN_0;
input 	Add5;
input 	Add51;
input 	in_ready_hold;
output 	in_data_reg_69;
output 	stateST_COMP_TRANS;
input 	mem_used_1;
output 	in_narrow_reg1;
input 	cp_ready;
output 	nxt_in_ready;
output 	out_valid_reg1;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready1;
input 	altera_reset_synchronizer_int_chain_out;
input 	Decoder1;
input 	Add2;
input 	Add21;
input 	Add22;
input 	Add23;
output 	nxt_in_ready2;
input 	src_valid;
output 	nxt_out_eop;
output 	out_byte_cnt_reg_2;
input 	cp_ready1;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_6;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_4;
output 	in_data_reg_105;
output 	in_data_reg_106;
output 	in_data_reg_107;
output 	in_data_reg_108;
output 	in_data_reg_109;
output 	in_data_reg_110;
output 	in_data_reg_111;
output 	in_data_reg_112;
output 	in_data_reg_113;
output 	in_data_reg_114;
output 	in_data_reg_115;
output 	in_data_reg_116;
input 	Selector10;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
input 	nxt_out_burstwrap_1;
input 	nxt_addr_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \align_address_to_size|LessThan0~0_combout ;
wire \align_address_to_size|LessThan0~1_combout ;
wire \NON_PIPELINED_INPUTS.load_next_cmd~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt[3]~1_combout ;
wire \Add4~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt[6]~2_combout ;
wire \nxt_uncomp_subburst_byte_cnt[5]~3_combout ;
wire \nxt_uncomp_subburst_byte_cnt[4]~4_combout ;
wire \nxt_uncomp_subburst_byte_cnt[2]~5_combout ;
wire \WideNor1~combout ;
wire \Selector2~1_combout ;
wire \load_next_out_cmd~combout ;
wire \state.ST_UNCOMP_TRANS~q ;
wire \Selector2~0_combout ;
wire \Selector0~0_combout ;
wire \state.ST_IDLE~q ;
wire \Selector1~0_combout ;
wire \Selector1~1_combout ;
wire \int_bytes_remaining_reg[4]~q ;
wire \d0_int_bytes_remaining[2]~1_combout ;
wire \int_bytes_remaining_reg[2]~q ;
wire \d0_int_bytes_remaining[3]~2_combout ;
wire \int_bytes_remaining_reg[3]~q ;
wire \Add1~0_combout ;
wire \d0_int_bytes_remaining[4]~0_combout ;
wire \int_bytes_remaining_reg[5]~q ;
wire \Add1~1_combout ;
wire \d0_int_bytes_remaining[5]~3_combout ;
wire \int_bytes_remaining_reg[6]~q ;
wire \d0_int_bytes_remaining[6]~4_combout ;
wire \new_burst_reg~0_combout ;
wire \new_burst_reg~q ;
wire \in_bytecount_reg_zero~0_combout ;
wire \in_bytecount_reg_zero~q ;
wire \nxt_out_valid~0_combout ;
wire \nxt_out_valid~1_combout ;
wire \Selector3~0_combout ;
wire \in_burstwrap_reg[3]~q ;
wire \nxt_addr[3]~0_combout ;
wire \nxt_addr[3]~combout ;
wire \int_nxt_addr_reg[3]~q ;
wire \in_size_reg[0]~q ;
wire \in_size_reg[1]~q ;
wire \in_size_reg[2]~q ;
wire \ShiftLeft0~0_combout ;
wire \ShiftLeft0~1_combout ;
wire \int_byte_cnt_narrow_reg[3]~q ;
wire \ShiftLeft0~2_combout ;
wire \int_byte_cnt_narrow_reg[2]~q ;
wire \in_burstwrap_reg[1]~q ;
wire \nxt_addr[1]~combout ;
wire \int_nxt_addr_reg[1]~q ;
wire \ShiftLeft0~3_combout ;
wire \int_byte_cnt_narrow_reg[1]~q ;
wire \int_byte_cnt_narrow_reg[0]~q ;
wire \Add0~13_sumout ;
wire \in_burstwrap_reg[0]~q ;
wire \nxt_addr[0]~combout ;
wire \int_nxt_addr_reg[0]~q ;
wire \d0_int_nxt_addr[0]~2_combout ;
wire \d0_int_nxt_addr[0]~3_combout ;
wire \int_nxt_addr_reg_dly[0]~q ;
wire \Add0~14 ;
wire \Add0~9_sumout ;
wire \d0_int_nxt_addr[1]~4_combout ;
wire \int_nxt_addr_reg_dly[1]~q ;
wire \Add0~10 ;
wire \Add0~6 ;
wire \Add0~1_sumout ;
wire \d0_int_nxt_addr[3]~0_combout ;
wire \in_burstwrap_reg[2]~q ;
wire \nxt_addr[2]~1_combout ;
wire \nxt_addr[2]~combout ;
wire \int_nxt_addr_reg[2]~q ;
wire \Add0~5_sumout ;
wire \d0_int_nxt_addr[2]~1_combout ;


spw_babasu_altera_merlin_address_alignment_16 align_address_to_size(
	.new_burst_reg(\new_burst_reg~q ),
	.src_payload(sink0_data[86]),
	.in_size_reg_0(\in_size_reg[0]~q ),
	.src_payload1(sink0_data[87]),
	.in_size_reg_1(\in_size_reg[1]~q ),
	.src_payload2(sink0_data[88]),
	.in_size_reg_2(\in_size_reg[2]~q ),
	.LessThan0(\align_address_to_size|LessThan0~0_combout ),
	.LessThan01(\align_address_to_size|LessThan0~1_combout ));

dffeas \in_data_reg[69] (
	.clk(clk_clk),
	.d(sink0_data[69]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_69),
	.prn(vcc));
defparam \in_data_reg[69] .is_wysiwyg = "true";
defparam \in_data_reg[69] .power_up = "low";

dffeas \state.ST_COMP_TRANS (
	.clk(clk_clk),
	.d(\Selector1~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_COMP_TRANS),
	.prn(vcc));
defparam \state.ST_COMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_COMP_TRANS .power_up = "low";

dffeas in_narrow_reg(
	.clk(clk_clk),
	.d(Decoder1),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_narrow_reg1),
	.prn(vcc));
defparam in_narrow_reg.is_wysiwyg = "true";
defparam in_narrow_reg.power_up = "low";

cyclonev_lcell_comb \nxt_in_ready~0 (
	.dataa(gnd),
	.datab(!stateST_COMP_TRANS),
	.datac(!\new_burst_reg~q ),
	.datad(!mem_used_1),
	.datae(!cp_ready),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~0 .extended_lut = "off";
defparam \nxt_in_ready~0 .lut_mask = 64'h0000030000000300;
defparam \nxt_in_ready~0 .shared_arith = "off";

dffeas out_valid_reg(
	.clk(clk_clk),
	.d(\nxt_out_valid~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_valid_reg1),
	.prn(vcc));
defparam out_valid_reg.is_wysiwyg = "true";
defparam out_valid_reg.power_up = "low";

dffeas \state.ST_UNCOMP_WR_SUBBURST (
	.clk(clk_clk),
	.d(\Selector3~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_UNCOMP_WR_SUBBURST),
	.prn(vcc));
defparam \state.ST_UNCOMP_WR_SUBBURST .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_WR_SUBBURST .power_up = "low";

cyclonev_lcell_comb \nxt_in_ready~1 (
	.dataa(!in_ready_hold),
	.datab(!stateST_COMP_TRANS),
	.datac(!mem_used_1),
	.datad(!cp_ready),
	.datae(!out_valid_reg1),
	.dataf(!\Selector2~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~1 .extended_lut = "off";
defparam \nxt_in_ready~1 .lut_mask = 64'h0000FF3F8888BBBB;
defparam \nxt_in_ready~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_in_ready~2 (
	.dataa(!nxt_in_ready),
	.datab(!nxt_in_ready1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready2),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~2 .extended_lut = "off";
defparam \nxt_in_ready~2 .lut_mask = 64'h2222222222222222;
defparam \nxt_in_ready~2 .shared_arith = "off";

cyclonev_lcell_comb \nxt_out_eop~0 (
	.dataa(!in_data_reg_69),
	.datab(!stateST_COMP_TRANS),
	.datac(!\new_burst_reg~q ),
	.datad(!mem_used_1),
	.datae(!cp_ready),
	.dataf(!\in_bytecount_reg_zero~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_out_eop),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_eop~0 .extended_lut = "off";
defparam \nxt_out_eop~0 .lut_mask = 64'h4444474477774777;
defparam \nxt_out_eop~0 .shared_arith = "off";

dffeas \out_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[3] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[3]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_3),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[3] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[3] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[2]~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[6] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[6]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_6),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[6] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[6] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[5] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[5]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_5),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[5] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[5] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[4] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[4]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_4),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[4] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[4] .power_up = "low";

dffeas \in_data_reg[105] (
	.clk(clk_clk),
	.d(sink0_data[105]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_105),
	.prn(vcc));
defparam \in_data_reg[105] .is_wysiwyg = "true";
defparam \in_data_reg[105] .power_up = "low";

dffeas \in_data_reg[106] (
	.clk(clk_clk),
	.d(sink0_data[106]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_106),
	.prn(vcc));
defparam \in_data_reg[106] .is_wysiwyg = "true";
defparam \in_data_reg[106] .power_up = "low";

dffeas \in_data_reg[107] (
	.clk(clk_clk),
	.d(sink0_data[107]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_107),
	.prn(vcc));
defparam \in_data_reg[107] .is_wysiwyg = "true";
defparam \in_data_reg[107] .power_up = "low";

dffeas \in_data_reg[108] (
	.clk(clk_clk),
	.d(sink0_data[108]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_108),
	.prn(vcc));
defparam \in_data_reg[108] .is_wysiwyg = "true";
defparam \in_data_reg[108] .power_up = "low";

dffeas \in_data_reg[109] (
	.clk(clk_clk),
	.d(sink0_data[109]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_109),
	.prn(vcc));
defparam \in_data_reg[109] .is_wysiwyg = "true";
defparam \in_data_reg[109] .power_up = "low";

dffeas \in_data_reg[110] (
	.clk(clk_clk),
	.d(sink0_data[110]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_110),
	.prn(vcc));
defparam \in_data_reg[110] .is_wysiwyg = "true";
defparam \in_data_reg[110] .power_up = "low";

dffeas \in_data_reg[111] (
	.clk(clk_clk),
	.d(sink0_data[111]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_111),
	.prn(vcc));
defparam \in_data_reg[111] .is_wysiwyg = "true";
defparam \in_data_reg[111] .power_up = "low";

dffeas \in_data_reg[112] (
	.clk(clk_clk),
	.d(sink0_data[112]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_112),
	.prn(vcc));
defparam \in_data_reg[112] .is_wysiwyg = "true";
defparam \in_data_reg[112] .power_up = "low";

dffeas \in_data_reg[113] (
	.clk(clk_clk),
	.d(sink0_data[113]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_113),
	.prn(vcc));
defparam \in_data_reg[113] .is_wysiwyg = "true";
defparam \in_data_reg[113] .power_up = "low";

dffeas \in_data_reg[114] (
	.clk(clk_clk),
	.d(sink0_data[114]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_114),
	.prn(vcc));
defparam \in_data_reg[114] .is_wysiwyg = "true";
defparam \in_data_reg[114] .power_up = "low";

dffeas \in_data_reg[115] (
	.clk(clk_clk),
	.d(sink0_data[115]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_115),
	.prn(vcc));
defparam \in_data_reg[115] .is_wysiwyg = "true";
defparam \in_data_reg[115] .power_up = "low";

dffeas \in_data_reg[116] (
	.clk(clk_clk),
	.d(sink0_data[116]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_116),
	.prn(vcc));
defparam \in_data_reg[116] .is_wysiwyg = "true";
defparam \in_data_reg[116] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[3] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[3]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_3),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[3] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[2] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[2]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_2),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[2] .power_up = "low";

cyclonev_lcell_comb \NON_PIPELINED_INPUTS.load_next_cmd~0 (
	.dataa(!in_ready_hold),
	.datab(!nxt_in_ready2),
	.datac(!src_valid),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \NON_PIPELINED_INPUTS.load_next_cmd~0 .extended_lut = "off";
defparam \NON_PIPELINED_INPUTS.load_next_cmd~0 .lut_mask = 64'h0404040404040404;
defparam \NON_PIPELINED_INPUTS.load_next_cmd~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt~0 (
	.dataa(!mem_used_1),
	.datab(!cp_ready),
	.datac(!out_valid_reg1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt~0 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt~0 .lut_mask = 64'h0202020202020202;
defparam \nxt_uncomp_subburst_byte_cnt~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[3]~1 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!out_uncomp_byte_cnt_reg_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[3]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[3]~1 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[3]~1 .lut_mask = 64'h0FE40F4E0FE40F4E;
defparam \nxt_uncomp_subburst_byte_cnt[3]~1 .shared_arith = "off";

cyclonev_lcell_comb \Add4~0 (
	.dataa(!out_uncomp_byte_cnt_reg_3),
	.datab(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datac(!out_uncomp_byte_cnt_reg_2),
	.datad(!out_uncomp_byte_cnt_reg_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add4~0 .extended_lut = "off";
defparam \Add4~0 .lut_mask = 64'h2000200020002000;
defparam \Add4~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[6]~2 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_6),
	.datae(!out_uncomp_byte_cnt_reg_5),
	.dataf(!\Add4~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[6]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[6]~2 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[6]~2 .lut_mask = 64'h04FE04FEAE5404FE;
defparam \nxt_uncomp_subburst_byte_cnt[6]~2 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[5]~3 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_5),
	.datae(!\Add4~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[5]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[5]~3 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[5]~3 .lut_mask = 64'h04FEAE5404FEAE54;
defparam \nxt_uncomp_subburst_byte_cnt[5]~3 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[4]~4 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!out_uncomp_byte_cnt_reg_2),
	.dataf(!out_uncomp_byte_cnt_reg_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[4]~4 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[4]~4 .lut_mask = 64'h00E40044FF4EFFEE;
defparam \nxt_uncomp_subburst_byte_cnt[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[2]~5 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[2]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[2]~5 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[2]~5 .lut_mask = 64'h0EF40EF40EF40EF4;
defparam \nxt_uncomp_subburst_byte_cnt[2]~5 .shared_arith = "off";

cyclonev_lcell_comb WideNor1(
	.dataa(!\nxt_uncomp_subburst_byte_cnt[3]~1_combout ),
	.datab(!\nxt_uncomp_subburst_byte_cnt[6]~2_combout ),
	.datac(!\nxt_uncomp_subburst_byte_cnt[5]~3_combout ),
	.datad(!\nxt_uncomp_subburst_byte_cnt[4]~4_combout ),
	.datae(!\nxt_uncomp_subburst_byte_cnt[2]~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideNor1.extended_lut = "off";
defparam WideNor1.lut_mask = 64'h8000000080000000;
defparam WideNor1.shared_arith = "off";

cyclonev_lcell_comb \Selector2~1 (
	.dataa(!nxt_out_eop),
	.datab(!\Selector2~0_combout ),
	.datac(!\WideNor1~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~1 .extended_lut = "off";
defparam \Selector2~1 .lut_mask = 64'h0808080808080808;
defparam \Selector2~1 .shared_arith = "off";

cyclonev_lcell_comb load_next_out_cmd(
	.dataa(!mem_used_1),
	.datab(!cp_ready),
	.datac(!out_valid_reg1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\load_next_out_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam load_next_out_cmd.extended_lut = "off";
defparam load_next_out_cmd.lut_mask = 64'hF2F2F2F2F2F2F2F2;
defparam load_next_out_cmd.shared_arith = "off";

dffeas \state.ST_UNCOMP_TRANS (
	.clk(clk_clk),
	.d(\Selector2~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_UNCOMP_TRANS~q ),
	.prn(vcc));
defparam \state.ST_UNCOMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_TRANS .power_up = "low";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'h8888888888888888;
defparam \Selector2~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!in_ready_hold),
	.datab(!nxt_out_eop),
	.datac(!src_valid),
	.datad(!\state.ST_IDLE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'h05CD05CD05CD05CD;
defparam \Selector0~0 .shared_arith = "off";

dffeas \state.ST_IDLE (
	.clk(clk_clk),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_IDLE~q ),
	.prn(vcc));
defparam \state.ST_IDLE .is_wysiwyg = "true";
defparam \state.ST_IDLE .power_up = "low";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!sink0_data[69]),
	.datab(!nxt_out_eop),
	.datac(!\Selector2~0_combout ),
	.datad(!\state.ST_IDLE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'h5510551055105510;
defparam \Selector1~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~1 (
	.dataa(!in_ready_hold),
	.datab(!stateST_COMP_TRANS),
	.datac(!nxt_out_eop),
	.datad(!src_valid),
	.datae(!\Selector1~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~1 .extended_lut = "off";
defparam \Selector1~1 .lut_mask = 64'h3031307530313075;
defparam \Selector1~1 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[4] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[4]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[4]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[4] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[4] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[2]~1 (
	.dataa(!h2f_ARLEN_0),
	.datab(!sink0_data[69]),
	.datac(!\new_burst_reg~q ),
	.datad(!out_byte_cnt_reg_2),
	.datae(!\int_bytes_remaining_reg[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[2]~1 .extended_lut = "off";
defparam \d0_int_bytes_remaining[2]~1 .lut_mask = 64'h02F2F20202F2F202;
defparam \d0_int_bytes_remaining[2]~1 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[2] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[2]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[2]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[2] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[3]~2 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!Add2),
	.datad(!\int_bytes_remaining_reg[3]~q ),
	.datae(!out_byte_cnt_reg_2),
	.dataf(!\int_bytes_remaining_reg[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[3]~2 .extended_lut = "off";
defparam \d0_int_bytes_remaining[3]~2 .lut_mask = 64'h01CDCD0101CD01CD;
defparam \d0_int_bytes_remaining[3]~2 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[3] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[3]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[3]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[3] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[3] .power_up = "low";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!\int_bytes_remaining_reg[4]~q ),
	.datab(!\int_bytes_remaining_reg[3]~q ),
	.datac(!out_byte_cnt_reg_2),
	.datad(!\int_bytes_remaining_reg[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'hA6AAA6AAA6AAA6AA;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[4]~0 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!Add21),
	.datad(!\Add1~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[4]~0 .extended_lut = "off";
defparam \d0_int_bytes_remaining[4]~0 .lut_mask = 64'hCD01CD01CD01CD01;
defparam \d0_int_bytes_remaining[4]~0 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[5] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[5]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[5]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[5] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[5] .power_up = "low";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!\int_bytes_remaining_reg[4]~q ),
	.datab(!\int_bytes_remaining_reg[3]~q ),
	.datac(!out_byte_cnt_reg_2),
	.datad(!\int_bytes_remaining_reg[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h0800080008000800;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[5]~3 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!Add22),
	.datad(!\int_bytes_remaining_reg[5]~q ),
	.datae(!\Add1~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[5]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[5]~3 .extended_lut = "off";
defparam \d0_int_bytes_remaining[5]~3 .lut_mask = 64'h01CDCD0101CDCD01;
defparam \d0_int_bytes_remaining[5]~3 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[6] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[6]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[6]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[6] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[6] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[6]~4 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!Add23),
	.datad(!\int_bytes_remaining_reg[5]~q ),
	.datae(!\Add1~1_combout ),
	.dataf(!\int_bytes_remaining_reg[6]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[6]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[6]~4 .extended_lut = "off";
defparam \d0_int_bytes_remaining[6]~4 .lut_mask = 64'h0101CD01CDCD01CD;
defparam \d0_int_bytes_remaining[6]~4 .shared_arith = "off";

cyclonev_lcell_comb \new_burst_reg~0 (
	.dataa(!\Selector1~1_combout ),
	.datab(!\d0_int_bytes_remaining[4]~0_combout ),
	.datac(!\d0_int_bytes_remaining[2]~1_combout ),
	.datad(!\d0_int_bytes_remaining[3]~2_combout ),
	.datae(!\d0_int_bytes_remaining[5]~3_combout ),
	.dataf(!\d0_int_bytes_remaining[6]~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\new_burst_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \new_burst_reg~0 .extended_lut = "off";
defparam \new_burst_reg~0 .lut_mask = 64'hAEAAAAAAAAAAAAAA;
defparam \new_burst_reg~0 .shared_arith = "off";

dffeas new_burst_reg(
	.clk(clk_clk),
	.d(\new_burst_reg~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\new_burst_reg~q ),
	.prn(vcc));
defparam new_burst_reg.is_wysiwyg = "true";
defparam new_burst_reg.power_up = "low";

cyclonev_lcell_comb \in_bytecount_reg_zero~0 (
	.dataa(!sink0_data[69]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\in_bytecount_reg_zero~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \in_bytecount_reg_zero~0 .extended_lut = "off";
defparam \in_bytecount_reg_zero~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \in_bytecount_reg_zero~0 .shared_arith = "off";

dffeas in_bytecount_reg_zero(
	.clk(clk_clk),
	.d(\in_bytecount_reg_zero~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_bytecount_reg_zero~q ),
	.prn(vcc));
defparam in_bytecount_reg_zero.is_wysiwyg = "true";
defparam in_bytecount_reg_zero.power_up = "low";

cyclonev_lcell_comb \nxt_out_valid~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!mem_used_1),
	.datac(!\in_bytecount_reg_zero~q ),
	.datad(!cp_ready1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_valid~0 .extended_lut = "off";
defparam \nxt_out_valid~0 .lut_mask = 64'hF0B8F0B8F0B8F0B8;
defparam \nxt_out_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_out_valid~1 (
	.dataa(!in_ready_hold),
	.datab(!stateST_COMP_TRANS),
	.datac(!src_valid),
	.datad(!\nxt_out_valid~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_valid~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_valid~1 .extended_lut = "off";
defparam \nxt_out_valid~1 .lut_mask = 64'h0537053705370537;
defparam \nxt_out_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~0 (
	.dataa(!nxt_out_eop),
	.datab(!\Selector2~0_combout ),
	.datac(!\WideNor1~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'h8080808080808080;
defparam \Selector3~0 .shared_arith = "off";

dffeas \in_burstwrap_reg[3] (
	.clk(clk_clk),
	.d(sink0_data[82]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_burstwrap_reg[3]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[3] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[3] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[3]~0 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!\in_burstwrap_reg[3]~q ),
	.datad(!\d0_int_nxt_addr[3]~0_combout ),
	.datae(!h2f_ARBURST_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[3]~0 .extended_lut = "off";
defparam \nxt_addr[3]~0 .lut_mask = 64'h00F300E200F300E2;
defparam \nxt_addr[3]~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_addr[3] (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!h2f_ARBURST_1),
	.datad(!Add5),
	.datae(!Selector10),
	.dataf(!\nxt_addr[3]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[3] .extended_lut = "off";
defparam \nxt_addr[3] .lut_mask = 64'h00000000FEEEFFEF;
defparam \nxt_addr[3] .shared_arith = "off";

dffeas \int_nxt_addr_reg[3] (
	.clk(clk_clk),
	.d(\nxt_addr[3]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[3]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[3] .power_up = "low";

dffeas \in_size_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[86]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_size_reg[0]~q ),
	.prn(vcc));
defparam \in_size_reg[0] .is_wysiwyg = "true";
defparam \in_size_reg[0] .power_up = "low";

dffeas \in_size_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[87]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_size_reg[1]~q ),
	.prn(vcc));
defparam \in_size_reg[1] .is_wysiwyg = "true";
defparam \in_size_reg[1] .power_up = "low";

dffeas \in_size_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[88]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_size_reg[2]~q ),
	.prn(vcc));
defparam \in_size_reg[2] .is_wysiwyg = "true";
defparam \in_size_reg[2] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[87]),
	.datac(!\in_size_reg[1]~q ),
	.datad(!sink0_data[88]),
	.datae(!\in_size_reg[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~0 .extended_lut = "off";
defparam \ShiftLeft0~0 .lut_mask = 64'h1B0A11001B0A1100;
defparam \ShiftLeft0~0 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~1 .extended_lut = "off";
defparam \ShiftLeft0~1 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~1 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[3] (
	.clk(clk_clk),
	.d(\ShiftLeft0~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[3]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[3] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[3] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~2 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~2 .extended_lut = "off";
defparam \ShiftLeft0~2 .lut_mask = 64'h00E400E400E400E4;
defparam \ShiftLeft0~2 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[2] (
	.clk(clk_clk),
	.d(\ShiftLeft0~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[2]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[2] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[2] .power_up = "low";

dffeas \in_burstwrap_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[80]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_burstwrap_reg[1]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[1] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[1] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[1] (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!\in_burstwrap_reg[1]~q ),
	.datad(!\d0_int_nxt_addr[1]~4_combout ),
	.datae(!nxt_out_burstwrap_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[1] .extended_lut = "off";
defparam \nxt_addr[1] .lut_mask = 64'h00E200F300E200F3;
defparam \nxt_addr[1] .shared_arith = "off";

dffeas \int_nxt_addr_reg[1] (
	.clk(clk_clk),
	.d(\nxt_addr[1]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[1] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\align_address_to_size|LessThan0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~3 .extended_lut = "off";
defparam \ShiftLeft0~3 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~3 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[1] (
	.clk(clk_clk),
	.d(\ShiftLeft0~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[1]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[1] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[1] .power_up = "low";

dffeas \int_byte_cnt_narrow_reg[0] (
	.clk(clk_clk),
	.d(\align_address_to_size|LessThan0~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[0]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[0] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[0] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[0]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \in_burstwrap_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[79]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_burstwrap_reg[0]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[0] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[0] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[0] (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!sink0_data[79]),
	.datad(!\in_burstwrap_reg[0]~q ),
	.datae(!\d0_int_nxt_addr[0]~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[0] .extended_lut = "off";
defparam \nxt_addr[0] .lut_mask = 64'h0000FE320000FE32;
defparam \nxt_addr[0] .shared_arith = "off";

dffeas \int_nxt_addr_reg[0] (
	.clk(clk_clk),
	.d(\nxt_addr[0]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[0] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~2 (
	.dataa(!\Add0~13_sumout ),
	.datab(!\int_nxt_addr_reg[0]~q ),
	.datac(!\in_burstwrap_reg[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~2 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~2 .lut_mask = 64'hC8C8C8C8C8C8C8C8;
defparam \d0_int_nxt_addr[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~3 (
	.dataa(!h2f_ARADDR_0),
	.datab(!sink0_data[69]),
	.datac(!\new_burst_reg~q ),
	.datad(!\align_address_to_size|LessThan0~1_combout ),
	.datae(!\d0_int_nxt_addr[0]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~3 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~3 .lut_mask = 64'hF0F10001F0F10001;
defparam \d0_int_nxt_addr[0]~3 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[0] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[0]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[0] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[1]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[1]~q ),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~4 (
	.dataa(!\int_nxt_addr_reg[1]~q ),
	.datab(!\Add0~9_sumout ),
	.datac(!sink0_data[69]),
	.datad(!Decoder1),
	.datae(!\new_burst_reg~q ),
	.dataf(!h2f_ARADDR_1),
	.datag(!\in_burstwrap_reg[1]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~4 .extended_lut = "on";
defparam \d0_int_nxt_addr[1]~4 .lut_mask = 64'h575700005757000F;
defparam \d0_int_nxt_addr[1]~4 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[1] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[1]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[1] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_2),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[2]~q ),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[3]~q ),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~0 (
	.dataa(!h2f_ARADDR_3),
	.datab(!sink0_data[69]),
	.datac(!\new_burst_reg~q ),
	.datad(!\int_nxt_addr_reg[3]~q ),
	.datae(!\in_burstwrap_reg[3]~q ),
	.dataf(!\Add0~1_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~0 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~0 .lut_mask = 64'h01F101F101F1F1F1;
defparam \d0_int_nxt_addr[3]~0 .shared_arith = "off";

dffeas \in_burstwrap_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[81]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_burstwrap_reg[2]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[2] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[2] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[2]~1 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!\in_burstwrap_reg[2]~q ),
	.datad(!\d0_int_nxt_addr[2]~1_combout ),
	.datae(!h2f_ARBURST_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[2]~1 .extended_lut = "off";
defparam \nxt_addr[2]~1 .lut_mask = 64'h00F300E200F300E2;
defparam \nxt_addr[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_addr[2] (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!h2f_ARBURST_1),
	.datad(!Add51),
	.datae(!\nxt_addr[2]~1_combout ),
	.dataf(!nxt_addr_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[2] .extended_lut = "off";
defparam \nxt_addr[2] .lut_mask = 64'h0000FEEE0000FFEF;
defparam \nxt_addr[2] .shared_arith = "off";

dffeas \int_nxt_addr_reg[2] (
	.clk(clk_clk),
	.d(\nxt_addr[2]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[2]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~1 (
	.dataa(!h2f_ARADDR_2),
	.datab(!sink0_data[69]),
	.datac(!\new_burst_reg~q ),
	.datad(!\int_nxt_addr_reg[2]~q ),
	.datae(!\in_burstwrap_reg[2]~q ),
	.dataf(!\Add0~5_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~1 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~1 .lut_mask = 64'h01F101F101F1F1F1;
defparam \d0_int_nxt_addr[2]~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_address_alignment_16 (
	new_burst_reg,
	src_payload,
	in_size_reg_0,
	src_payload1,
	in_size_reg_1,
	src_payload2,
	in_size_reg_2,
	LessThan0,
	LessThan01)/* synthesis synthesis_greybox=0 */;
input 	new_burst_reg;
input 	src_payload;
input 	in_size_reg_0;
input 	src_payload1;
input 	in_size_reg_1;
input 	src_payload2;
input 	in_size_reg_2;
output 	LessThan0;
output 	LessThan01;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!new_burst_reg),
	.datab(!src_payload1),
	.datac(!in_size_reg_1),
	.datad(!src_payload2),
	.datae(!in_size_reg_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan0),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'hE4A04400E4A04400;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~1 (
	.dataa(!new_burst_reg),
	.datab(!src_payload),
	.datac(!in_size_reg_0),
	.datad(!LessThan0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan01),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~1 .extended_lut = "off";
defparam \LessThan0~1 .lut_mask = 64'h00E400E400E400E4;
defparam \LessThan0~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_burst_adapter_16 (
	h2f_ARADDR_0,
	h2f_ARADDR_1,
	h2f_ARADDR_2,
	h2f_ARADDR_3,
	h2f_ARLEN_0,
	nxt_in_ready,
	in_ready_hold,
	stateST_COMP_TRANS,
	out_valid_reg,
	in_narrow_reg,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	in_data_reg_68,
	cp_ready,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready1,
	saved_grant_1,
	Equal5,
	saved_grant_0,
	altera_reset_synchronizer_int_chain_out,
	in_data_reg_0,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	Add2,
	Add21,
	Add22,
	Add23,
	write_cp_data_77,
	write_cp_data_78,
	write_cp_data_75,
	write_cp_data_74,
	write_cp_data_76,
	WideNor0,
	Equal14,
	nxt_out_eop,
	src6_valid,
	src_valid,
	cp_ready1,
	in_data_reg_69,
	src_data_87,
	src_data_88,
	src_valid1,
	src_data_35,
	src_data_34,
	src_data_33,
	src_data_32,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_6,
	src_payload_0,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	Selector3,
	Selector10,
	base_address_3,
	Selector4,
	Selector11,
	base_address_2,
	src_payload,
	src_data_82,
	src_data_81,
	src_data_105,
	src_data_106,
	src_data_107,
	src_data_108,
	src_data_109,
	src_data_110,
	src_data_111,
	src_data_112,
	src_data_113,
	src_data_114,
	src_data_115,
	src_data_116,
	src_data_86,
	Selector5,
	Selector12,
	out_data_1,
	src_data_80,
	out_data_0,
	Selector6,
	Selector13,
	src_data_79,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARADDR_0;
input 	h2f_ARADDR_1;
input 	h2f_ARADDR_2;
input 	h2f_ARADDR_3;
input 	h2f_ARLEN_0;
output 	nxt_in_ready;
input 	in_ready_hold;
output 	stateST_COMP_TRANS;
output 	out_valid_reg;
output 	in_narrow_reg;
output 	in_byteen_reg_3;
output 	in_byteen_reg_2;
output 	in_byteen_reg_1;
output 	in_byteen_reg_0;
output 	in_data_reg_68;
input 	cp_ready;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready1;
input 	saved_grant_1;
input 	Equal5;
input 	saved_grant_0;
input 	altera_reset_synchronizer_int_chain_out;
output 	in_data_reg_0;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
input 	Add2;
input 	Add21;
input 	Add22;
input 	Add23;
input 	write_cp_data_77;
input 	write_cp_data_78;
input 	write_cp_data_75;
input 	write_cp_data_74;
input 	write_cp_data_76;
input 	WideNor0;
input 	Equal14;
output 	nxt_out_eop;
input 	src6_valid;
input 	src_valid;
input 	cp_ready1;
output 	in_data_reg_69;
input 	src_data_87;
input 	src_data_88;
input 	src_valid1;
input 	src_data_35;
input 	src_data_34;
input 	src_data_33;
input 	src_data_32;
output 	out_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_6;
input 	src_payload_0;
output 	in_data_reg_105;
output 	in_data_reg_106;
output 	in_data_reg_107;
output 	in_data_reg_108;
output 	in_data_reg_109;
output 	in_data_reg_110;
output 	in_data_reg_111;
output 	in_data_reg_112;
output 	in_data_reg_113;
output 	in_data_reg_114;
output 	in_data_reg_115;
output 	in_data_reg_116;
input 	Selector3;
input 	Selector10;
input 	base_address_3;
input 	Selector4;
input 	Selector11;
input 	base_address_2;
input 	src_payload;
input 	src_data_82;
input 	src_data_81;
input 	src_data_105;
input 	src_data_106;
input 	src_data_107;
input 	src_data_108;
input 	src_data_109;
input 	src_data_110;
input 	src_data_111;
input 	src_data_112;
input 	src_data_113;
input 	src_data_114;
input 	src_data_115;
input 	src_data_116;
input 	src_data_86;
input 	Selector5;
input 	Selector12;
input 	out_data_1;
input 	src_data_80;
input 	out_data_0;
input 	Selector6;
input 	Selector13;
input 	src_data_79;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



spw_babasu_altera_merlin_burst_adapter_13_1_16 \altera_merlin_burst_adapter_13_1.burst_adapter (
	.h2f_ARADDR_0(h2f_ARADDR_0),
	.h2f_ARADDR_1(h2f_ARADDR_1),
	.h2f_ARADDR_2(h2f_ARADDR_2),
	.h2f_ARADDR_3(h2f_ARADDR_3),
	.h2f_ARLEN_0(h2f_ARLEN_0),
	.nxt_in_ready(nxt_in_ready),
	.in_ready_hold(in_ready_hold),
	.stateST_COMP_TRANS(stateST_COMP_TRANS),
	.out_valid_reg1(out_valid_reg),
	.in_narrow_reg1(in_narrow_reg),
	.in_byteen_reg_3(in_byteen_reg_3),
	.in_byteen_reg_2(in_byteen_reg_2),
	.in_byteen_reg_1(in_byteen_reg_1),
	.in_byteen_reg_0(in_byteen_reg_0),
	.in_data_reg_68(in_data_reg_68),
	.cp_ready(cp_ready),
	.stateST_UNCOMP_WR_SUBBURST(stateST_UNCOMP_WR_SUBBURST),
	.nxt_in_ready1(nxt_in_ready1),
	.sink0_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_116,src_data_115,src_data_114,src_data_113,src_data_112,src_data_111,src_data_110,src_data_109,src_data_108,src_data_107,src_data_106,src_data_105,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_88,src_data_87,
src_data_86,gnd,gnd,gnd,src_data_82,src_data_81,src_data_80,src_data_79,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,saved_grant_1,saved_grant_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_35,src_data_34,src_data_33,
src_data_32,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_payload}),
	.Equal5(Equal5),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.in_data_reg_0(in_data_reg_0),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_3),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_2),
	.Add2(Add2),
	.Add21(Add21),
	.Add22(Add22),
	.Add23(Add23),
	.write_cp_data_77(write_cp_data_77),
	.write_cp_data_78(write_cp_data_78),
	.write_cp_data_75(write_cp_data_75),
	.write_cp_data_74(write_cp_data_74),
	.write_cp_data_76(write_cp_data_76),
	.WideNor0(WideNor0),
	.Equal14(Equal14),
	.nxt_out_eop(nxt_out_eop),
	.src6_valid(src6_valid),
	.src_valid(src_valid),
	.cp_ready1(cp_ready1),
	.in_data_reg_69(in_data_reg_69),
	.src_valid1(src_valid1),
	.out_byte_cnt_reg_2(out_byte_cnt_reg_2),
	.out_uncomp_byte_cnt_reg_4(out_uncomp_byte_cnt_reg_4),
	.out_uncomp_byte_cnt_reg_3(out_uncomp_byte_cnt_reg_3),
	.out_uncomp_byte_cnt_reg_2(out_uncomp_byte_cnt_reg_2),
	.out_uncomp_byte_cnt_reg_5(out_uncomp_byte_cnt_reg_5),
	.out_uncomp_byte_cnt_reg_6(out_uncomp_byte_cnt_reg_6),
	.sink0_endofpacket(src_payload_0),
	.in_data_reg_105(in_data_reg_105),
	.in_data_reg_106(in_data_reg_106),
	.in_data_reg_107(in_data_reg_107),
	.in_data_reg_108(in_data_reg_108),
	.in_data_reg_109(in_data_reg_109),
	.in_data_reg_110(in_data_reg_110),
	.in_data_reg_111(in_data_reg_111),
	.in_data_reg_112(in_data_reg_112),
	.in_data_reg_113(in_data_reg_113),
	.in_data_reg_114(in_data_reg_114),
	.in_data_reg_115(in_data_reg_115),
	.in_data_reg_116(in_data_reg_116),
	.Selector3(Selector3),
	.Selector10(Selector10),
	.base_address_3(base_address_3),
	.Selector4(Selector4),
	.Selector11(Selector11),
	.base_address_2(base_address_2),
	.Selector5(Selector5),
	.Selector12(Selector12),
	.out_data_1(out_data_1),
	.out_data_0(out_data_0),
	.Selector6(Selector6),
	.Selector13(Selector13),
	.clk_clk(clk_clk));

endmodule

module spw_babasu_altera_merlin_burst_adapter_13_1_16 (
	h2f_ARADDR_0,
	h2f_ARADDR_1,
	h2f_ARADDR_2,
	h2f_ARADDR_3,
	h2f_ARLEN_0,
	nxt_in_ready,
	in_ready_hold,
	stateST_COMP_TRANS,
	out_valid_reg1,
	in_narrow_reg1,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	in_data_reg_68,
	cp_ready,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready1,
	sink0_data,
	Equal5,
	altera_reset_synchronizer_int_chain_out,
	in_data_reg_0,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	Add2,
	Add21,
	Add22,
	Add23,
	write_cp_data_77,
	write_cp_data_78,
	write_cp_data_75,
	write_cp_data_74,
	write_cp_data_76,
	WideNor0,
	Equal14,
	nxt_out_eop,
	src6_valid,
	src_valid,
	cp_ready1,
	in_data_reg_69,
	src_valid1,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_6,
	sink0_endofpacket,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	in_data_reg_113,
	in_data_reg_114,
	in_data_reg_115,
	in_data_reg_116,
	Selector3,
	Selector10,
	base_address_3,
	Selector4,
	Selector11,
	base_address_2,
	Selector5,
	Selector12,
	out_data_1,
	out_data_0,
	Selector6,
	Selector13,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARADDR_0;
input 	h2f_ARADDR_1;
input 	h2f_ARADDR_2;
input 	h2f_ARADDR_3;
input 	h2f_ARLEN_0;
output 	nxt_in_ready;
input 	in_ready_hold;
output 	stateST_COMP_TRANS;
output 	out_valid_reg1;
output 	in_narrow_reg1;
output 	in_byteen_reg_3;
output 	in_byteen_reg_2;
output 	in_byteen_reg_1;
output 	in_byteen_reg_0;
output 	in_data_reg_68;
input 	cp_ready;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready1;
input 	[128:0] sink0_data;
input 	Equal5;
input 	altera_reset_synchronizer_int_chain_out;
output 	in_data_reg_0;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
input 	Add2;
input 	Add21;
input 	Add22;
input 	Add23;
input 	write_cp_data_77;
input 	write_cp_data_78;
input 	write_cp_data_75;
input 	write_cp_data_74;
input 	write_cp_data_76;
input 	WideNor0;
input 	Equal14;
output 	nxt_out_eop;
input 	src6_valid;
input 	src_valid;
input 	cp_ready1;
output 	in_data_reg_69;
input 	src_valid1;
output 	out_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_6;
input 	sink0_endofpacket;
output 	in_data_reg_105;
output 	in_data_reg_106;
output 	in_data_reg_107;
output 	in_data_reg_108;
output 	in_data_reg_109;
output 	in_data_reg_110;
output 	in_data_reg_111;
output 	in_data_reg_112;
output 	in_data_reg_113;
output 	in_data_reg_114;
output 	in_data_reg_115;
output 	in_data_reg_116;
input 	Selector3;
input 	Selector10;
input 	base_address_3;
input 	Selector4;
input 	Selector11;
input 	base_address_2;
input 	Selector5;
input 	Selector12;
input 	out_data_1;
input 	out_data_0;
input 	Selector6;
input 	Selector13;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \align_address_to_size|LessThan0~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt[4]~1_combout ;
wire \nxt_uncomp_subburst_byte_cnt[3]~2_combout ;
wire \Add4~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt[5]~3_combout ;
wire \nxt_uncomp_subburst_byte_cnt[2]~4_combout ;
wire \nxt_uncomp_subburst_byte_cnt[6]~5_combout ;
wire \WideOr0~combout ;
wire \in_valid~combout ;
wire \Selector0~0_combout ;
wire \load_next_out_cmd~combout ;
wire \state.ST_IDLE~q ;
wire \Selector2~0_combout ;
wire \Selector2~1_combout ;
wire \Selector2~2_combout ;
wire \state.ST_UNCOMP_TRANS~q ;
wire \Selector1~0_combout ;
wire \Selector1~1_combout ;
wire \int_bytes_remaining_reg[5]~q ;
wire \d0_int_bytes_remaining[2]~5_combout ;
wire \d0_int_bytes_remaining[2]~6_combout ;
wire \int_bytes_remaining_reg[2]~q ;
wire \d0_int_bytes_remaining[3]~7_combout ;
wire \d0_int_bytes_remaining[3]~8_combout ;
wire \int_bytes_remaining_reg[3]~q ;
wire \Add1~1_combout ;
wire \d0_int_bytes_remaining[4]~4_combout ;
wire \int_bytes_remaining_reg[4]~q ;
wire \Add1~0_combout ;
wire \d0_int_bytes_remaining[5]~0_combout ;
wire \d0_int_bytes_remaining[5]~1_combout ;
wire \int_bytes_remaining_reg[6]~q ;
wire \d0_int_bytes_remaining[6]~2_combout ;
wire \d0_int_bytes_remaining[6]~3_combout ;
wire \new_burst_reg~0_combout ;
wire \new_burst_reg~q ;
wire \WideNor0~0_combout ;
wire \NON_PIPELINED_INPUTS.load_next_cmd~combout ;
wire \in_bytecount_reg_zero~q ;
wire \nxt_out_valid~0_combout ;
wire \LessThan0~0_combout ;
wire \Selector3~0_combout ;
wire \in_size_reg[0]~q ;
wire \in_size_reg[2]~q ;
wire \in_size_reg[1]~q ;
wire \ShiftLeft0~0_combout ;
wire \ShiftLeft0~1_combout ;
wire \int_byte_cnt_narrow_reg[3]~q ;
wire \ShiftLeft0~2_combout ;
wire \int_byte_cnt_narrow_reg[2]~q ;
wire \ShiftLeft0~3_combout ;
wire \ShiftLeft0~4_combout ;
wire \int_byte_cnt_narrow_reg[1]~q ;
wire \int_byte_cnt_narrow_reg[0]~q ;
wire \Add0~13_sumout ;
wire \d0_int_nxt_addr[0]~3_combout ;
wire \in_burstwrap_reg[0]~q ;
wire \nxt_addr[0]~0_combout ;
wire \int_nxt_addr_reg[0]~q ;
wire \d0_int_nxt_addr[0]~4_combout ;
wire \int_nxt_addr_reg_dly[0]~q ;
wire \Add0~14 ;
wire \Add0~9_sumout ;
wire \in_burstwrap_reg[1]~q ;
wire \nxt_addr[1]~4_combout ;
wire \int_nxt_addr_reg[1]~q ;
wire \d0_int_nxt_addr[1]~7_combout ;
wire \d0_int_nxt_addr[1]~2_combout ;
wire \int_nxt_addr_reg_dly[1]~q ;
wire \Add0~10 ;
wire \Add0~6 ;
wire \Add0~1_sumout ;
wire \in_burstwrap_reg[3]~q ;
wire \nxt_addr[3]~12_combout ;
wire \int_nxt_addr_reg[3]~q ;
wire \d0_int_nxt_addr[3]~5_combout ;
wire \d0_int_nxt_addr[3]~0_combout ;
wire \Add0~5_sumout ;
wire \in_burstwrap_reg[2]~q ;
wire \nxt_addr[2]~8_combout ;
wire \int_nxt_addr_reg[2]~q ;
wire \d0_int_nxt_addr[2]~6_combout ;
wire \d0_int_nxt_addr[2]~1_combout ;
wire \in_eop_reg~q ;


spw_babasu_altera_merlin_address_alignment_17 align_address_to_size(
	.new_burst_reg(\new_burst_reg~q ),
	.src_data_86(sink0_data[86]),
	.in_size_reg_0(\in_size_reg[0]~q ),
	.ShiftLeft0(\ShiftLeft0~3_combout ),
	.LessThan0(\align_address_to_size|LessThan0~0_combout ));

cyclonev_lcell_comb \nxt_in_ready~1 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!in_ready_hold),
	.datac(!out_valid_reg1),
	.datad(!cp_ready),
	.datae(!stateST_COMP_TRANS),
	.dataf(!\new_burst_reg~q ),
	.datag(!stateST_UNCOMP_WR_SUBBURST),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~1 .extended_lut = "on";
defparam \nxt_in_ready~1 .lut_mask = 64'h2020F0F02020F0FF;
defparam \nxt_in_ready~1 .shared_arith = "off";

dffeas \state.ST_COMP_TRANS (
	.clk(clk_clk),
	.d(\Selector1~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_COMP_TRANS),
	.prn(vcc));
defparam \state.ST_COMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_COMP_TRANS .power_up = "low";

dffeas out_valid_reg(
	.clk(clk_clk),
	.d(\nxt_out_valid~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_valid_reg1),
	.prn(vcc));
defparam out_valid_reg.is_wysiwyg = "true";
defparam out_valid_reg.power_up = "low";

dffeas in_narrow_reg(
	.clk(clk_clk),
	.d(\LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_narrow_reg1),
	.prn(vcc));
defparam in_narrow_reg.is_wysiwyg = "true";
defparam in_narrow_reg.power_up = "low";

dffeas \in_byteen_reg[3] (
	.clk(clk_clk),
	.d(sink0_data[35]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_3),
	.prn(vcc));
defparam \in_byteen_reg[3] .is_wysiwyg = "true";
defparam \in_byteen_reg[3] .power_up = "low";

dffeas \in_byteen_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[34]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_2),
	.prn(vcc));
defparam \in_byteen_reg[2] .is_wysiwyg = "true";
defparam \in_byteen_reg[2] .power_up = "low";

dffeas \in_byteen_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[33]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_1),
	.prn(vcc));
defparam \in_byteen_reg[1] .is_wysiwyg = "true";
defparam \in_byteen_reg[1] .power_up = "low";

dffeas \in_byteen_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[32]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_0),
	.prn(vcc));
defparam \in_byteen_reg[0] .is_wysiwyg = "true";
defparam \in_byteen_reg[0] .power_up = "low";

dffeas \in_data_reg[68] (
	.clk(clk_clk),
	.d(sink0_data[68]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_68),
	.prn(vcc));
defparam \in_data_reg[68] .is_wysiwyg = "true";
defparam \in_data_reg[68] .power_up = "low";

dffeas \state.ST_UNCOMP_WR_SUBBURST (
	.clk(clk_clk),
	.d(\Selector3~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_UNCOMP_WR_SUBBURST),
	.prn(vcc));
defparam \state.ST_UNCOMP_WR_SUBBURST .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_WR_SUBBURST .power_up = "low";

cyclonev_lcell_comb \nxt_in_ready~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!out_valid_reg1),
	.datac(!cp_ready),
	.datad(!\state.ST_UNCOMP_TRANS~q ),
	.datae(!stateST_UNCOMP_WR_SUBBURST),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~0 .extended_lut = "off";
defparam \nxt_in_ready~0 .lut_mask = 64'h008A8A8A008A8A8A;
defparam \nxt_in_ready~0 .shared_arith = "off";

dffeas \in_data_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[0]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_0),
	.prn(vcc));
defparam \in_data_reg[0] .is_wysiwyg = "true";
defparam \in_data_reg[0] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[3] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[3]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_3),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[3] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[2] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[2]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_2),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[2] .power_up = "low";

cyclonev_lcell_comb \nxt_out_eop~0 (
	.dataa(!\in_eop_reg~q ),
	.datab(!stateST_COMP_TRANS),
	.datac(!\new_burst_reg~q ),
	.datad(!cp_ready),
	.datae(!\in_bytecount_reg_zero~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_out_eop),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_eop~0 .extended_lut = "off";
defparam \nxt_out_eop~0 .lut_mask = 64'h4447774744477747;
defparam \nxt_out_eop~0 .shared_arith = "off";

dffeas \in_data_reg[69] (
	.clk(clk_clk),
	.d(sink0_data[69]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_69),
	.prn(vcc));
defparam \in_data_reg[69] .is_wysiwyg = "true";
defparam \in_data_reg[69] .power_up = "low";

dffeas \out_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[4] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[4]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_4),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[4] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[4] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[3] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[3]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_3),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[3] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[3] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[2]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[5] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[5]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_5),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[5] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[5] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[6] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[6]~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_6),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[6] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[6] .power_up = "low";

dffeas \in_data_reg[105] (
	.clk(clk_clk),
	.d(sink0_data[105]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_105),
	.prn(vcc));
defparam \in_data_reg[105] .is_wysiwyg = "true";
defparam \in_data_reg[105] .power_up = "low";

dffeas \in_data_reg[106] (
	.clk(clk_clk),
	.d(sink0_data[106]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_106),
	.prn(vcc));
defparam \in_data_reg[106] .is_wysiwyg = "true";
defparam \in_data_reg[106] .power_up = "low";

dffeas \in_data_reg[107] (
	.clk(clk_clk),
	.d(sink0_data[107]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_107),
	.prn(vcc));
defparam \in_data_reg[107] .is_wysiwyg = "true";
defparam \in_data_reg[107] .power_up = "low";

dffeas \in_data_reg[108] (
	.clk(clk_clk),
	.d(sink0_data[108]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_108),
	.prn(vcc));
defparam \in_data_reg[108] .is_wysiwyg = "true";
defparam \in_data_reg[108] .power_up = "low";

dffeas \in_data_reg[109] (
	.clk(clk_clk),
	.d(sink0_data[109]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_109),
	.prn(vcc));
defparam \in_data_reg[109] .is_wysiwyg = "true";
defparam \in_data_reg[109] .power_up = "low";

dffeas \in_data_reg[110] (
	.clk(clk_clk),
	.d(sink0_data[110]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_110),
	.prn(vcc));
defparam \in_data_reg[110] .is_wysiwyg = "true";
defparam \in_data_reg[110] .power_up = "low";

dffeas \in_data_reg[111] (
	.clk(clk_clk),
	.d(sink0_data[111]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_111),
	.prn(vcc));
defparam \in_data_reg[111] .is_wysiwyg = "true";
defparam \in_data_reg[111] .power_up = "low";

dffeas \in_data_reg[112] (
	.clk(clk_clk),
	.d(sink0_data[112]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_112),
	.prn(vcc));
defparam \in_data_reg[112] .is_wysiwyg = "true";
defparam \in_data_reg[112] .power_up = "low";

dffeas \in_data_reg[113] (
	.clk(clk_clk),
	.d(sink0_data[113]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_113),
	.prn(vcc));
defparam \in_data_reg[113] .is_wysiwyg = "true";
defparam \in_data_reg[113] .power_up = "low";

dffeas \in_data_reg[114] (
	.clk(clk_clk),
	.d(sink0_data[114]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_114),
	.prn(vcc));
defparam \in_data_reg[114] .is_wysiwyg = "true";
defparam \in_data_reg[114] .power_up = "low";

dffeas \in_data_reg[115] (
	.clk(clk_clk),
	.d(sink0_data[115]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_115),
	.prn(vcc));
defparam \in_data_reg[115] .is_wysiwyg = "true";
defparam \in_data_reg[115] .power_up = "low";

dffeas \in_data_reg[116] (
	.clk(clk_clk),
	.d(sink0_data[116]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_116),
	.prn(vcc));
defparam \in_data_reg[116] .is_wysiwyg = "true";
defparam \in_data_reg[116] .power_up = "low";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt~0 (
	.dataa(!out_valid_reg1),
	.datab(!cp_ready),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt~0 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt~0 .lut_mask = 64'h1111111111111111;
defparam \nxt_uncomp_subburst_byte_cnt~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[4]~1 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!out_uncomp_byte_cnt_reg_3),
	.datae(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.dataf(!out_uncomp_byte_cnt_reg_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[4]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[4]~1 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[4]~1 .lut_mask = 64'h0F0FE44E0F0F4E4E;
defparam \nxt_uncomp_subburst_byte_cnt[4]~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[3]~2 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!out_uncomp_byte_cnt_reg_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[3]~2 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[3]~2 .lut_mask = 64'h0FE40F4E0FE40F4E;
defparam \nxt_uncomp_subburst_byte_cnt[3]~2 .shared_arith = "off";

cyclonev_lcell_comb \Add4~0 (
	.dataa(!out_uncomp_byte_cnt_reg_4),
	.datab(!out_uncomp_byte_cnt_reg_3),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add4~0 .extended_lut = "off";
defparam \Add4~0 .lut_mask = 64'h0800080008000800;
defparam \Add4~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[5]~3 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_5),
	.datae(!\Add4~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[5]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[5]~3 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[5]~3 .lut_mask = 64'h04FEAE5404FEAE54;
defparam \nxt_uncomp_subburst_byte_cnt[5]~3 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[2]~4 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[2]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[2]~4 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[2]~4 .lut_mask = 64'h0EF40EF40EF40EF4;
defparam \nxt_uncomp_subburst_byte_cnt[2]~4 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[6]~5 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_5),
	.datae(!\Add4~0_combout ),
	.dataf(!out_uncomp_byte_cnt_reg_6),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[6]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[6]~5 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[6]~5 .lut_mask = 64'h0404AE04FEFE54FE;
defparam \nxt_uncomp_subburst_byte_cnt[6]~5 .shared_arith = "off";

cyclonev_lcell_comb WideOr0(
	.dataa(!\nxt_uncomp_subburst_byte_cnt[4]~1_combout ),
	.datab(!\nxt_uncomp_subburst_byte_cnt[3]~2_combout ),
	.datac(!\nxt_uncomp_subburst_byte_cnt[5]~3_combout ),
	.datad(!\nxt_uncomp_subburst_byte_cnt[2]~4_combout ),
	.datae(!\nxt_uncomp_subburst_byte_cnt[6]~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr0.extended_lut = "off";
defparam WideOr0.lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam WideOr0.shared_arith = "off";

cyclonev_lcell_comb in_valid(
	.dataa(!in_ready_hold),
	.datab(!Equal5),
	.datac(!Equal14),
	.datad(!sink0_data[68]),
	.datae(!src6_valid),
	.dataf(!src_valid),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\in_valid~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam in_valid.extended_lut = "off";
defparam in_valid.lut_mask = 64'h0000000155555555;
defparam in_valid.shared_arith = "off";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!sink0_data[69]),
	.datab(!nxt_out_eop),
	.datac(!sink0_data[68]),
	.datad(!\in_valid~combout ),
	.datae(!\state.ST_IDLE~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'h005FCCFF005FCCFF;
defparam \Selector0~0 .shared_arith = "off";

cyclonev_lcell_comb load_next_out_cmd(
	.dataa(!out_valid_reg1),
	.datab(!cp_ready),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\load_next_out_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam load_next_out_cmd.extended_lut = "off";
defparam load_next_out_cmd.lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam load_next_out_cmd.shared_arith = "off";

dffeas \state.ST_IDLE (
	.clk(clk_clk),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_IDLE~q ),
	.prn(vcc));
defparam \state.ST_IDLE .is_wysiwyg = "true";
defparam \state.ST_IDLE .power_up = "low";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!nxt_out_eop),
	.datac(!stateST_UNCOMP_WR_SUBBURST),
	.datad(!\state.ST_IDLE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'h00EC00EC00EC00EC;
defparam \Selector2~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~1 (
	.dataa(!in_ready_hold),
	.datab(!Equal5),
	.datac(!Equal14),
	.datad(!sink0_data[68]),
	.datae(!src6_valid),
	.dataf(!\Selector2~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~1 .extended_lut = "off";
defparam \Selector2~1 .lut_mask = 64'h0000000100000000;
defparam \Selector2~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~2 (
	.dataa(!\WideOr0~combout ),
	.datab(!\Selector2~1_combout ),
	.datac(!\in_valid~combout ),
	.datad(!nxt_out_eop),
	.datae(!\state.ST_UNCOMP_TRANS~q ),
	.dataf(!sink0_data[69]),
	.datag(!stateST_UNCOMP_WR_SUBBURST),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~2 .extended_lut = "on";
defparam \Selector2~2 .lut_mask = 64'h3B33BB3F0A00AA00;
defparam \Selector2~2 .shared_arith = "off";

dffeas \state.ST_UNCOMP_TRANS (
	.clk(clk_clk),
	.d(\Selector2~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_UNCOMP_TRANS~q ),
	.prn(vcc));
defparam \state.ST_UNCOMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_TRANS .power_up = "low";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!nxt_out_eop),
	.datac(!\state.ST_UNCOMP_TRANS~q ),
	.datad(!stateST_UNCOMP_WR_SUBBURST),
	.datae(!\state.ST_IDLE~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'h0000A8880000A888;
defparam \Selector1~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~1 (
	.dataa(!sink0_data[69]),
	.datab(!stateST_COMP_TRANS),
	.datac(!nxt_out_eop),
	.datad(!sink0_data[68]),
	.datae(!\in_valid~combout ),
	.dataf(!\Selector1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~1 .extended_lut = "off";
defparam \Selector1~1 .lut_mask = 64'h3030777530303330;
defparam \Selector1~1 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[5] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[5]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[5]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[5] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[5] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[2]~5 (
	.dataa(!h2f_ARLEN_0),
	.datab(!sink0_data[69]),
	.datac(!sink0_data[68]),
	.datad(!write_cp_data_74),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[2]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[2]~5 .extended_lut = "off";
defparam \d0_int_bytes_remaining[2]~5 .lut_mask = 64'h2F222F222F222F22;
defparam \d0_int_bytes_remaining[2]~5 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[2]~6 (
	.dataa(!\new_burst_reg~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\int_bytes_remaining_reg[2]~q ),
	.datad(!\d0_int_bytes_remaining[2]~5_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[2]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[2]~6 .extended_lut = "off";
defparam \d0_int_bytes_remaining[2]~6 .lut_mask = 64'h287D287D287D287D;
defparam \d0_int_bytes_remaining[2]~6 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[2] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[2]~6_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[2]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[2] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[3]~7 (
	.dataa(!sink0_data[69]),
	.datab(!sink0_data[68]),
	.datac(!write_cp_data_75),
	.datad(!Add2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[3]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[3]~7 .extended_lut = "off";
defparam \d0_int_bytes_remaining[3]~7 .lut_mask = 64'h0357035703570357;
defparam \d0_int_bytes_remaining[3]~7 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[3]~8 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\int_bytes_remaining_reg[3]~q ),
	.datac(!out_byte_cnt_reg_2),
	.datad(!\int_bytes_remaining_reg[2]~q ),
	.datae(!\d0_int_bytes_remaining[3]~7_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[3]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[3]~8 .extended_lut = "off";
defparam \d0_int_bytes_remaining[3]~8 .lut_mask = 64'h28227D7728227D77;
defparam \d0_int_bytes_remaining[3]~8 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[3] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[3]~8_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[3]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[3] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[3] .power_up = "low";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!\int_bytes_remaining_reg[4]~q ),
	.datab(!\int_bytes_remaining_reg[3]~q ),
	.datac(!out_byte_cnt_reg_2),
	.datad(!\int_bytes_remaining_reg[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'hA6AAA6AAA6AAA6AA;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[4]~4 (
	.dataa(!sink0_data[69]),
	.datab(!\new_burst_reg~q ),
	.datac(!sink0_data[68]),
	.datad(!write_cp_data_76),
	.datae(!Add21),
	.dataf(!\Add1~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[4]~4 .extended_lut = "off";
defparam \d0_int_bytes_remaining[4]~4 .lut_mask = 64'hCCCFDDDF00031113;
defparam \d0_int_bytes_remaining[4]~4 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[4] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[4]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[4]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[4] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[4] .power_up = "low";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!\int_bytes_remaining_reg[4]~q ),
	.datab(!\int_bytes_remaining_reg[3]~q ),
	.datac(!out_byte_cnt_reg_2),
	.datad(!\int_bytes_remaining_reg[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h0800080008000800;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[5]~0 (
	.dataa(!sink0_data[69]),
	.datab(!sink0_data[68]),
	.datac(!write_cp_data_77),
	.datad(!Add22),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[5]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[5]~0 .extended_lut = "off";
defparam \d0_int_bytes_remaining[5]~0 .lut_mask = 64'h0357035703570357;
defparam \d0_int_bytes_remaining[5]~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[5]~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\int_bytes_remaining_reg[5]~q ),
	.datac(!\Add1~0_combout ),
	.datad(!\d0_int_bytes_remaining[5]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[5]~1 .extended_lut = "off";
defparam \d0_int_bytes_remaining[5]~1 .lut_mask = 64'h287D287D287D287D;
defparam \d0_int_bytes_remaining[5]~1 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[6] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[6]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[6]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[6] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[6] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[6]~2 (
	.dataa(!sink0_data[69]),
	.datab(!sink0_data[68]),
	.datac(!write_cp_data_78),
	.datad(!Add23),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[6]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[6]~2 .extended_lut = "off";
defparam \d0_int_bytes_remaining[6]~2 .lut_mask = 64'h0357035703570357;
defparam \d0_int_bytes_remaining[6]~2 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[6]~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\int_bytes_remaining_reg[5]~q ),
	.datac(!\Add1~0_combout ),
	.datad(!\int_bytes_remaining_reg[6]~q ),
	.datae(!\d0_int_bytes_remaining[6]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[6]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[6]~3 .extended_lut = "off";
defparam \d0_int_bytes_remaining[6]~3 .lut_mask = 64'h08A25DF708A25DF7;
defparam \d0_int_bytes_remaining[6]~3 .shared_arith = "off";

cyclonev_lcell_comb \new_burst_reg~0 (
	.dataa(!\Selector1~1_combout ),
	.datab(!\d0_int_bytes_remaining[5]~1_combout ),
	.datac(!\d0_int_bytes_remaining[6]~3_combout ),
	.datad(!\d0_int_bytes_remaining[4]~4_combout ),
	.datae(!\d0_int_bytes_remaining[2]~6_combout ),
	.dataf(!\d0_int_bytes_remaining[3]~8_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\new_burst_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \new_burst_reg~0 .extended_lut = "off";
defparam \new_burst_reg~0 .lut_mask = 64'hAAAAEAAAAAAAAAAA;
defparam \new_burst_reg~0 .shared_arith = "off";

dffeas new_burst_reg(
	.clk(clk_clk),
	.d(\new_burst_reg~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\new_burst_reg~q ),
	.prn(vcc));
defparam new_burst_reg.is_wysiwyg = "true";
defparam new_burst_reg.power_up = "low";

cyclonev_lcell_comb \WideNor0~0 (
	.dataa(!sink0_data[69]),
	.datab(!sink0_data[68]),
	.datac(!WideNor0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideNor0~0 .extended_lut = "off";
defparam \WideNor0~0 .lut_mask = 64'h8A8A8A8A8A8A8A8A;
defparam \WideNor0~0 .shared_arith = "off";

cyclonev_lcell_comb \NON_PIPELINED_INPUTS.load_next_cmd (
	.dataa(!in_ready_hold),
	.datab(!nxt_in_ready1),
	.datac(!nxt_in_ready),
	.datad(!src_valid),
	.datae(!src_valid1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \NON_PIPELINED_INPUTS.load_next_cmd .extended_lut = "off";
defparam \NON_PIPELINED_INPUTS.load_next_cmd .lut_mask = 64'h0015151500151515;
defparam \NON_PIPELINED_INPUTS.load_next_cmd .shared_arith = "off";

dffeas in_bytecount_reg_zero(
	.clk(clk_clk),
	.d(\WideNor0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_bytecount_reg_zero~q ),
	.prn(vcc));
defparam in_bytecount_reg_zero.is_wysiwyg = "true";
defparam in_bytecount_reg_zero.power_up = "low";

cyclonev_lcell_comb \nxt_out_valid~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!\new_burst_reg~q ),
	.datac(!\in_bytecount_reg_zero~q ),
	.datad(!\in_valid~combout ),
	.datae(!cp_ready1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_valid~0 .extended_lut = "off";
defparam \nxt_out_valid~0 .lut_mask = 64'h50FF44FF50FF44FF;
defparam \nxt_out_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!sink0_data[87]),
	.datab(!sink0_data[88]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h8888888888888888;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~0 (
	.dataa(!nxt_out_eop),
	.datab(!\state.ST_UNCOMP_TRANS~q ),
	.datac(!stateST_UNCOMP_WR_SUBBURST),
	.datad(!\WideOr0~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'h002A002A002A002A;
defparam \Selector3~0 .shared_arith = "off";

dffeas \in_size_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[86]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[0]~q ),
	.prn(vcc));
defparam \in_size_reg[0] .is_wysiwyg = "true";
defparam \in_size_reg[0] .power_up = "low";

dffeas \in_size_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[88]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[2]~q ),
	.prn(vcc));
defparam \in_size_reg[2] .is_wysiwyg = "true";
defparam \in_size_reg[2] .power_up = "low";

dffeas \in_size_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[87]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[1]~q ),
	.prn(vcc));
defparam \in_size_reg[1] .is_wysiwyg = "true";
defparam \in_size_reg[1] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[87]),
	.datac(!sink0_data[88]),
	.datad(!\in_size_reg[2]~q ),
	.datae(!\in_size_reg[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~0 .extended_lut = "off";
defparam \ShiftLeft0~0 .lut_mask = 64'h1010BA101010BA10;
defparam \ShiftLeft0~0 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~1 .extended_lut = "off";
defparam \ShiftLeft0~1 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~1 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[3] (
	.clk(clk_clk),
	.d(\ShiftLeft0~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[3]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[3] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[3] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~2 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~2 .extended_lut = "off";
defparam \ShiftLeft0~2 .lut_mask = 64'h00E400E400E400E4;
defparam \ShiftLeft0~2 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[2] (
	.clk(clk_clk),
	.d(\ShiftLeft0~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[2]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[2] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[2] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[87]),
	.datac(!sink0_data[88]),
	.datad(!\in_size_reg[2]~q ),
	.datae(!\in_size_reg[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~3 .extended_lut = "off";
defparam \ShiftLeft0~3 .lut_mask = 64'hEA404040EA404040;
defparam \ShiftLeft0~3 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~4 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[86]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~4 .extended_lut = "off";
defparam \ShiftLeft0~4 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~4 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[1] (
	.clk(clk_clk),
	.d(\ShiftLeft0~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[1]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[1] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[1] .power_up = "low";

dffeas \int_byte_cnt_narrow_reg[0] (
	.clk(clk_clk),
	.d(\align_address_to_size|LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[0]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[0] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[0] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[0]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~3 (
	.dataa(!h2f_ARADDR_0),
	.datab(!sink0_data[69]),
	.datac(!sink0_data[68]),
	.datad(!out_data_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~3 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~3 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[0]~3 .shared_arith = "off";

dffeas \in_burstwrap_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[79]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[0]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[0] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[0] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[0]~0 (
	.dataa(!Selector13),
	.datab(!Selector6),
	.datac(!sink0_data[68]),
	.datad(!sink0_data[69]),
	.datae(!\new_burst_reg~q ),
	.dataf(!\d0_int_nxt_addr[0]~4_combout ),
	.datag(!\in_burstwrap_reg[0]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[0]~0 .extended_lut = "on";
defparam \nxt_addr[0]~0 .lut_mask = 64'h00000000F0F0FCA8;
defparam \nxt_addr[0]~0 .shared_arith = "off";

dffeas \int_nxt_addr_reg[0] (
	.clk(clk_clk),
	.d(\nxt_addr[0]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[0] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~4 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\Add0~13_sumout ),
	.datac(!\align_address_to_size|LessThan0~0_combout ),
	.datad(!\d0_int_nxt_addr[0]~3_combout ),
	.datae(!\int_nxt_addr_reg[0]~q ),
	.dataf(!\in_burstwrap_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~4 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~4 .lut_mask = 64'h0005AAAF2227AAAF;
defparam \d0_int_nxt_addr[0]~4 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[0] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[0]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[0] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[1]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[1]~q ),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \in_burstwrap_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[80]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[1]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[1] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[1] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[1]~4 (
	.dataa(!Selector12),
	.datab(!Selector5),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!\new_burst_reg~q ),
	.dataf(!\d0_int_nxt_addr[1]~2_combout ),
	.datag(!\in_burstwrap_reg[1]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[1]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[1]~4 .extended_lut = "on";
defparam \nxt_addr[1]~4 .lut_mask = 64'h00000000F0F0FAC8;
defparam \nxt_addr[1]~4 .shared_arith = "off";

dffeas \int_nxt_addr_reg[1] (
	.clk(clk_clk),
	.d(\nxt_addr[1]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[1] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~7 (
	.dataa(!h2f_ARADDR_1),
	.datab(!sink0_data[69]),
	.datac(!sink0_data[68]),
	.datad(!out_data_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~7 .extended_lut = "off";
defparam \d0_int_nxt_addr[1]~7 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[1]~7 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~2 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\Add0~9_sumout ),
	.datac(!\in_burstwrap_reg[1]~q ),
	.datad(!\int_nxt_addr_reg[1]~q ),
	.datae(!\ShiftLeft0~3_combout ),
	.dataf(!\d0_int_nxt_addr[1]~7_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~2 .extended_lut = "off";
defparam \d0_int_nxt_addr[1]~2 .lut_mask = 64'h02AA02AA02AA57FF;
defparam \d0_int_nxt_addr[1]~2 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[1] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[1]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[1] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_2),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[2]~q ),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[3]~q ),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

dffeas \in_burstwrap_reg[3] (
	.clk(clk_clk),
	.d(sink0_data[82]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[3]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[3] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[3] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[3]~12 (
	.dataa(!Selector10),
	.datab(!Selector3),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!\new_burst_reg~q ),
	.dataf(!\d0_int_nxt_addr[3]~0_combout ),
	.datag(!\in_burstwrap_reg[3]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[3]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[3]~12 .extended_lut = "on";
defparam \nxt_addr[3]~12 .lut_mask = 64'h00000000F0F0FAC8;
defparam \nxt_addr[3]~12 .shared_arith = "off";

dffeas \int_nxt_addr_reg[3] (
	.clk(clk_clk),
	.d(\nxt_addr[3]~12_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[3]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[3] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~5 (
	.dataa(!\Add0~1_sumout ),
	.datab(!\in_burstwrap_reg[3]~q ),
	.datac(!\int_nxt_addr_reg[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~5 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~5 .lut_mask = 64'hE0E0E0E0E0E0E0E0;
defparam \d0_int_nxt_addr[3]~5 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!h2f_ARADDR_3),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!base_address_3),
	.dataf(!\d0_int_nxt_addr[3]~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~0 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~0 .lut_mask = 64'hABABABFF01010155;
defparam \d0_int_nxt_addr[3]~0 .shared_arith = "off";

dffeas \in_burstwrap_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[81]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[2]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[2] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[2] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[2]~8 (
	.dataa(!Selector11),
	.datab(!Selector4),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!\new_burst_reg~q ),
	.dataf(!\d0_int_nxt_addr[2]~1_combout ),
	.datag(!\in_burstwrap_reg[2]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[2]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[2]~8 .extended_lut = "on";
defparam \nxt_addr[2]~8 .lut_mask = 64'h00000000F0F0FAC8;
defparam \nxt_addr[2]~8 .shared_arith = "off";

dffeas \int_nxt_addr_reg[2] (
	.clk(clk_clk),
	.d(\nxt_addr[2]~8_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[2]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~6 (
	.dataa(!\Add0~5_sumout ),
	.datab(!\in_burstwrap_reg[2]~q ),
	.datac(!\int_nxt_addr_reg[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~6 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~6 .lut_mask = 64'hE0E0E0E0E0E0E0E0;
defparam \d0_int_nxt_addr[2]~6 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!h2f_ARADDR_2),
	.datac(!sink0_data[69]),
	.datad(!sink0_data[68]),
	.datae(!base_address_2),
	.dataf(!\d0_int_nxt_addr[2]~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~1 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~1 .lut_mask = 64'hABABABFF01010155;
defparam \d0_int_nxt_addr[2]~1 .shared_arith = "off";

dffeas in_eop_reg(
	.clk(clk_clk),
	.d(sink0_endofpacket),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_eop_reg~q ),
	.prn(vcc));
defparam in_eop_reg.is_wysiwyg = "true";
defparam in_eop_reg.power_up = "low";

endmodule

module spw_babasu_altera_merlin_address_alignment_17 (
	new_burst_reg,
	src_data_86,
	in_size_reg_0,
	ShiftLeft0,
	LessThan0)/* synthesis synthesis_greybox=0 */;
input 	new_burst_reg;
input 	src_data_86;
input 	in_size_reg_0;
input 	ShiftLeft0;
output 	LessThan0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!new_burst_reg),
	.datab(!src_data_86),
	.datac(!in_size_reg_0),
	.datad(!ShiftLeft0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan0),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h00E400E400E400E4;
defparam \LessThan0~0 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_slave_agent (
	waitrequest_reset_override,
	stateST_COMP_TRANS,
	out_valid_reg,
	mem_used_1,
	in_narrow_reg,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	WideOr0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	in_data_reg_68,
	cp_ready,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_129_0,
	mem_used_01,
	mem_66_0,
	comb,
	last_packet_beat,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	last_packet_beat1,
	m0_write1,
	altera_reset_synchronizer_int_chain_out,
	nxt_out_eop,
	cp_ready1,
	last_packet_beat2,
	WideOr01,
	read,
	cp_ready2,
	in_data_reg_69,
	rf_source_valid,
	rf_sink_ready,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	waitrequest_reset_override;
input 	stateST_COMP_TRANS;
input 	out_valid_reg;
input 	mem_used_1;
input 	in_narrow_reg;
input 	in_byteen_reg_3;
input 	in_byteen_reg_2;
input 	in_byteen_reg_1;
input 	in_byteen_reg_0;
output 	WideOr0;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	in_data_reg_68;
output 	cp_ready;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	mem_129_0;
input 	mem_used_01;
input 	mem_66_0;
output 	comb;
output 	last_packet_beat;
input 	mem_78_0;
input 	mem_77_0;
input 	mem_76_0;
input 	mem_75_0;
input 	mem_74_0;
output 	last_packet_beat1;
output 	m0_write1;
input 	altera_reset_synchronizer_int_chain_out;
input 	nxt_out_eop;
output 	cp_ready1;
output 	last_packet_beat2;
input 	WideOr01;
input 	read;
output 	cp_ready2;
input 	in_data_reg_69;
output 	rf_source_valid;
output 	rf_sink_ready;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \local_write~combout ;
wire \cp_ready~1_combout ;
wire \cp_ready~2_combout ;


spw_babasu_altera_merlin_burst_uncompressor uncompressor(
	.mem_66_0(mem_66_0),
	.comb(comb),
	.last_packet_beat(last_packet_beat),
	.mem_78_0(mem_78_0),
	.mem_77_0(mem_77_0),
	.mem_76_0(mem_76_0),
	.mem_75_0(mem_75_0),
	.mem_74_0(mem_74_0),
	.last_packet_beat1(last_packet_beat1),
	.reset(altera_reset_synchronizer_int_chain_out),
	.last_packet_beat2(last_packet_beat2),
	.WideOr0(WideOr01),
	.read(read),
	.sink_ready(rf_sink_ready),
	.clk(clk_clk));

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!in_narrow_reg),
	.datac(!in_byteen_reg_3),
	.datad(!in_byteen_reg_2),
	.datae(!in_byteen_reg_1),
	.dataf(!in_byteen_reg_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h1FFFFFFFFFFFFFFF;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~0 (
	.dataa(!waitrequest_reset_override),
	.datab(!mem_used_1),
	.datac(!WideOr0),
	.datad(!wait_latency_counter_1),
	.datae(!wait_latency_counter_0),
	.dataf(!\local_write~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~0 .extended_lut = "off";
defparam \cp_ready~0 .lut_mask = 64'hC0C0C4C0C4C0C0C0;
defparam \cp_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \comb~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_129_0),
	.datad(!mem_used_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(comb),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~0 .extended_lut = "off";
defparam \comb~0 .lut_mask = 64'h007F007F007F007F;
defparam \comb~0 .shared_arith = "off";

cyclonev_lcell_comb m0_write(
	.dataa(!mem_used_1),
	.datab(!WideOr0),
	.datac(!\local_write~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write1),
	.sumout(),
	.cout(),
	.shareout());
defparam m0_write.extended_lut = "off";
defparam m0_write.lut_mask = 64'h0202020202020202;
defparam m0_write.shared_arith = "off";

cyclonev_lcell_comb \cp_ready~3 (
	.dataa(!mem_used_1),
	.datab(!in_narrow_reg),
	.datac(!\cp_ready~1_combout ),
	.datad(!\cp_ready~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~3 .extended_lut = "off";
defparam \cp_ready~3 .lut_mask = 64'h08AA08AA08AA08AA;
defparam \cp_ready~3 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~4 (
	.dataa(!waitrequest_reset_override),
	.datab(!mem_used_1),
	.datac(!WideOr0),
	.datad(!wait_latency_counter_1),
	.datae(!wait_latency_counter_0),
	.dataf(!\local_write~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready2),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~4 .extended_lut = "off";
defparam \cp_ready~4 .lut_mask = 64'h0000550004005100;
defparam \cp_ready~4 .shared_arith = "off";

cyclonev_lcell_comb \rf_source_valid~0 (
	.dataa(!in_data_reg_68),
	.datab(!out_valid_reg),
	.datac(!nxt_out_eop),
	.datad(!in_data_reg_69),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rf_source_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_source_valid~0 .extended_lut = "off";
defparam \rf_source_valid~0 .lut_mask = 64'h0133013301330133;
defparam \rf_source_valid~0 .shared_arith = "off";

cyclonev_lcell_comb local_write(
	.dataa(!in_data_reg_68),
	.datab(!out_valid_reg),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\local_write~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam local_write.extended_lut = "off";
defparam local_write.lut_mask = 64'h1111111111111111;
defparam local_write.shared_arith = "off";

cyclonev_lcell_comb \cp_ready~1 (
	.dataa(!in_byteen_reg_3),
	.datab(!in_byteen_reg_2),
	.datac(!in_byteen_reg_1),
	.datad(!in_byteen_reg_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cp_ready~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~1 .extended_lut = "off";
defparam \cp_ready~1 .lut_mask = 64'h8000800080008000;
defparam \cp_ready~1 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~2 (
	.dataa(!waitrequest_reset_override),
	.datab(!wait_latency_counter_1),
	.datac(!wait_latency_counter_0),
	.datad(!\local_write~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cp_ready~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~2 .extended_lut = "off";
defparam \cp_ready~2 .lut_mask = 64'h0440044004400440;
defparam \cp_ready~2 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_burst_uncompressor (
	mem_66_0,
	comb,
	last_packet_beat,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	last_packet_beat1,
	reset,
	last_packet_beat2,
	WideOr0,
	read,
	sink_ready,
	clk)/* synthesis synthesis_greybox=0 */;
input 	mem_66_0;
input 	comb;
output 	last_packet_beat;
input 	mem_78_0;
input 	mem_77_0;
input 	mem_76_0;
input 	mem_75_0;
input 	mem_74_0;
output 	last_packet_beat1;
input 	reset;
output 	last_packet_beat2;
input 	WideOr0;
input 	read;
output 	sink_ready;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \burst_uncompress_busy~q ;
wire \burst_uncompress_byte_counter~5_combout ;
wire \burst_uncompress_byte_counter[2]~q ;
wire \burst_uncompress_byte_counter~4_combout ;
wire \burst_uncompress_byte_counter[3]~q ;
wire \Add0~2_combout ;
wire \burst_uncompress_byte_counter~3_combout ;
wire \burst_uncompress_byte_counter[4]~q ;
wire \last_packet_beat~3_combout ;
wire \Add1~0_combout ;
wire \burst_uncompress_byte_counter~6_combout ;
wire \burst_uncompress_byte_counter[7]~q ;
wire \burst_uncompress_byte_counter~0_combout ;
wire \Add0~1_combout ;
wire \Add1~1_combout ;
wire \burst_uncompress_byte_counter~2_combout ;
wire \burst_uncompress_byte_counter[5]~q ;
wire \Add0~0_combout ;
wire \burst_uncompress_byte_counter~1_combout ;
wire \burst_uncompress_byte_counter[6]~q ;


cyclonev_lcell_comb \last_packet_beat~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!\burst_uncompress_byte_counter[5]~q ),
	.datad(!\burst_uncompress_byte_counter[4]~q ),
	.datae(!\burst_uncompress_byte_counter[3]~q ),
	.dataf(!\burst_uncompress_byte_counter[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~0 .extended_lut = "off";
defparam \last_packet_beat~0 .lut_mask = 64'h0000000040000000;
defparam \last_packet_beat~0 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~1 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_78_0),
	.datac(!mem_77_0),
	.datad(!mem_76_0),
	.datae(!mem_75_0),
	.dataf(!mem_74_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat1),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~1 .extended_lut = "off";
defparam \last_packet_beat~1 .lut_mask = 64'h0000000080000000;
defparam \last_packet_beat~1 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~2 (
	.dataa(!comb),
	.datab(!mem_66_0),
	.datac(!last_packet_beat),
	.datad(!last_packet_beat1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat2),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~2 .extended_lut = "off";
defparam \last_packet_beat~2 .lut_mask = 64'h3222322232223222;
defparam \last_packet_beat~2 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!comb),
	.datad(!last_packet_beat2),
	.datae(!WideOr0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~0 .extended_lut = "off";
defparam \sink_ready~0 .lut_mask = 64'h00000F0000000F00;
defparam \sink_ready~0 .shared_arith = "off";

dffeas burst_uncompress_busy(
	.clk(clk),
	.d(last_packet_beat2),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_busy~q ),
	.prn(vcc));
defparam burst_uncompress_busy.is_wysiwyg = "true";
defparam burst_uncompress_busy.power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~5 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_74_0),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(!last_packet_beat2),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~5 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~5 .lut_mask = 64'h00C800FA00C800FA;
defparam \burst_uncompress_byte_counter~5 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[2] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[2]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[2] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[2] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~4 (
	.dataa(!mem_75_0),
	.datab(!mem_74_0),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(!last_packet_beat2),
	.dataf(!\burst_uncompress_byte_counter~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~4 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~4 .lut_mask = 64'h000099990000F00F;
defparam \burst_uncompress_byte_counter~4 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[3] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[3]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[3] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[3] .power_up = "low";

cyclonev_lcell_comb \Add0~2 (
	.dataa(!\burst_uncompress_byte_counter[4]~q ),
	.datab(!\burst_uncompress_byte_counter[3]~q ),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~2 .extended_lut = "off";
defparam \Add0~2 .lut_mask = 64'h6A6A6A6A6A6A6A6A;
defparam \Add0~2 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~3 (
	.dataa(!mem_76_0),
	.datab(!mem_75_0),
	.datac(!mem_74_0),
	.datad(!last_packet_beat2),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add0~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~3 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~3 .lut_mask = 64'h009500FF00950000;
defparam \burst_uncompress_byte_counter~3 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[4] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[4]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[4] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[4] .power_up = "low";

cyclonev_lcell_comb \last_packet_beat~3 (
	.dataa(!\burst_uncompress_byte_counter[6]~q ),
	.datab(!\burst_uncompress_byte_counter[5]~q ),
	.datac(!\burst_uncompress_byte_counter[4]~q ),
	.datad(!\burst_uncompress_byte_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_packet_beat~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~3 .extended_lut = "off";
defparam \last_packet_beat~3 .lut_mask = 64'h8000800080008000;
defparam \last_packet_beat~3 .shared_arith = "off";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!mem_77_0),
	.datab(!mem_76_0),
	.datac(!mem_75_0),
	.datad(!mem_74_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h8000800080008000;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~6 (
	.dataa(!mem_78_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat2),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~6 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~6 .lut_mask = 64'h0000000C0A0A000C;
defparam \burst_uncompress_byte_counter~6 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[7] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[7]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[7] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[7] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[2]~q ),
	.datac(!\last_packet_beat~3_combout ),
	.datad(!\burst_uncompress_byte_counter[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~0 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~0 .lut_mask = 64'h5155515551555155;
defparam \burst_uncompress_byte_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!mem_77_0),
	.datab(!mem_76_0),
	.datac(!mem_75_0),
	.datad(!mem_74_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~2 (
	.dataa(!last_packet_beat2),
	.datab(!\burst_uncompress_byte_counter~0_combout ),
	.datac(!\Add0~1_combout ),
	.datad(!\Add1~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~2 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~2 .lut_mask = 64'h5410541054105410;
defparam \burst_uncompress_byte_counter~2 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[5] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[5]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[5] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[5] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h8000800080008000;
defparam \Add0~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~1 (
	.dataa(!mem_78_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat2),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~1 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~1 .lut_mask = 64'h0505030C0A0A030C;
defparam \burst_uncompress_byte_counter~1 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[6] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[6]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[6] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[6] .power_up = "low";

endmodule

module spw_babasu_altera_merlin_slave_agent_1 (
	h2f_RREADY_0,
	waitrequest_reset_override,
	stateST_COMP_TRANS,
	mem_used_1,
	in_data_reg_69,
	in_narrow_reg,
	wait_latency_counter_1,
	wait_latency_counter_0,
	cp_ready,
	cp_ready1,
	empty,
	mem_66_0,
	mem_used_0,
	last_packet_beat,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	last_packet_beat1,
	altera_reset_synchronizer_int_chain_out,
	last_packet_beat2,
	cp_ready2,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_RREADY_0;
input 	waitrequest_reset_override;
input 	stateST_COMP_TRANS;
input 	mem_used_1;
input 	in_data_reg_69;
input 	in_narrow_reg;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
output 	cp_ready;
output 	cp_ready1;
input 	empty;
input 	mem_66_0;
input 	mem_used_0;
output 	last_packet_beat;
input 	mem_78_0;
input 	mem_77_0;
input 	mem_76_0;
input 	mem_75_0;
input 	mem_74_0;
output 	last_packet_beat1;
input 	altera_reset_synchronizer_int_chain_out;
output 	last_packet_beat2;
output 	cp_ready2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



spw_babasu_altera_merlin_burst_uncompressor_1 uncompressor(
	.h2f_RREADY_0(h2f_RREADY_0),
	.empty(empty),
	.mem_66_0(mem_66_0),
	.mem_used_0(mem_used_0),
	.last_packet_beat(last_packet_beat),
	.mem_78_0(mem_78_0),
	.mem_77_0(mem_77_0),
	.mem_76_0(mem_76_0),
	.mem_75_0(mem_75_0),
	.mem_74_0(mem_74_0),
	.last_packet_beat1(last_packet_beat1),
	.reset(altera_reset_synchronizer_int_chain_out),
	.last_packet_beat2(last_packet_beat2),
	.clk(clk_clk));

cyclonev_lcell_comb \cp_ready~0 (
	.dataa(!waitrequest_reset_override),
	.datab(!in_data_reg_69),
	.datac(!stateST_COMP_TRANS),
	.datad(!in_narrow_reg),
	.datae(!wait_latency_counter_1),
	.dataf(!wait_latency_counter_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~0 .extended_lut = "off";
defparam \cp_ready~0 .lut_mask = 64'hCCC0CCC0DDD5CCC0;
defparam \cp_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~1 (
	.dataa(!mem_used_1),
	.datab(!cp_ready),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~1 .extended_lut = "off";
defparam \cp_ready~1 .lut_mask = 64'h2222222222222222;
defparam \cp_ready~1 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~2 (
	.dataa(!waitrequest_reset_override),
	.datab(!in_data_reg_69),
	.datac(!in_narrow_reg),
	.datad(!wait_latency_counter_1),
	.datae(!wait_latency_counter_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready2),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~2 .extended_lut = "off";
defparam \cp_ready~2 .lut_mask = 64'hC0C0D5C0C0C0D5C0;
defparam \cp_ready~2 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_burst_uncompressor_1 (
	h2f_RREADY_0,
	empty,
	mem_66_0,
	mem_used_0,
	last_packet_beat,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	last_packet_beat1,
	reset,
	last_packet_beat2,
	clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_RREADY_0;
input 	empty;
input 	mem_66_0;
input 	mem_used_0;
output 	last_packet_beat;
input 	mem_78_0;
input 	mem_77_0;
input 	mem_76_0;
input 	mem_75_0;
input 	mem_74_0;
output 	last_packet_beat1;
input 	reset;
output 	last_packet_beat2;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always0~0_combout ;
wire \burst_uncompress_busy~q ;
wire \burst_uncompress_byte_counter~5_combout ;
wire \burst_uncompress_byte_counter[2]~q ;
wire \burst_uncompress_byte_counter~4_combout ;
wire \burst_uncompress_byte_counter[3]~q ;
wire \Add0~2_combout ;
wire \burst_uncompress_byte_counter~3_combout ;
wire \burst_uncompress_byte_counter[4]~q ;
wire \last_packet_beat~3_combout ;
wire \Add1~0_combout ;
wire \burst_uncompress_byte_counter~6_combout ;
wire \burst_uncompress_byte_counter[7]~q ;
wire \burst_uncompress_byte_counter~0_combout ;
wire \Add0~1_combout ;
wire \Add1~1_combout ;
wire \burst_uncompress_byte_counter~2_combout ;
wire \burst_uncompress_byte_counter[5]~q ;
wire \Add0~0_combout ;
wire \burst_uncompress_byte_counter~1_combout ;
wire \burst_uncompress_byte_counter[6]~q ;


cyclonev_lcell_comb \last_packet_beat~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!\burst_uncompress_byte_counter[5]~q ),
	.datad(!\burst_uncompress_byte_counter[4]~q ),
	.datae(!\burst_uncompress_byte_counter[3]~q ),
	.dataf(!\burst_uncompress_byte_counter[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~0 .extended_lut = "off";
defparam \last_packet_beat~0 .lut_mask = 64'h0000000040000000;
defparam \last_packet_beat~0 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~1 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_78_0),
	.datac(!mem_77_0),
	.datad(!mem_76_0),
	.datae(!mem_75_0),
	.dataf(!mem_74_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat1),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~1 .extended_lut = "off";
defparam \last_packet_beat~1 .lut_mask = 64'h0000000080000000;
defparam \last_packet_beat~1 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~2 (
	.dataa(!empty),
	.datab(!mem_66_0),
	.datac(!mem_used_0),
	.datad(!last_packet_beat),
	.datae(!last_packet_beat1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat2),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~2 .extended_lut = "off";
defparam \last_packet_beat~2 .lut_mask = 64'h3331313133313131;
defparam \last_packet_beat~2 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!h2f_RREADY_0),
	.datab(!empty),
	.datac(!mem_used_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'h0404040404040404;
defparam \always0~0 .shared_arith = "off";

dffeas burst_uncompress_busy(
	.clk(clk),
	.d(last_packet_beat2),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_busy~q ),
	.prn(vcc));
defparam burst_uncompress_busy.is_wysiwyg = "true";
defparam burst_uncompress_busy.power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~5 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_74_0),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(!last_packet_beat2),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~5 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~5 .lut_mask = 64'h00C800FA00C800FA;
defparam \burst_uncompress_byte_counter~5 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[2] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[2]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[2] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[2] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~4 (
	.dataa(!mem_75_0),
	.datab(!mem_74_0),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(!last_packet_beat2),
	.dataf(!\burst_uncompress_byte_counter~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~4 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~4 .lut_mask = 64'h000099990000F00F;
defparam \burst_uncompress_byte_counter~4 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[3] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[3]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[3] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[3] .power_up = "low";

cyclonev_lcell_comb \Add0~2 (
	.dataa(!\burst_uncompress_byte_counter[4]~q ),
	.datab(!\burst_uncompress_byte_counter[3]~q ),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~2 .extended_lut = "off";
defparam \Add0~2 .lut_mask = 64'h6A6A6A6A6A6A6A6A;
defparam \Add0~2 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~3 (
	.dataa(!mem_76_0),
	.datab(!mem_75_0),
	.datac(!mem_74_0),
	.datad(!last_packet_beat2),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add0~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~3 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~3 .lut_mask = 64'h009500FF00950000;
defparam \burst_uncompress_byte_counter~3 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[4] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[4]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[4] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[4] .power_up = "low";

cyclonev_lcell_comb \last_packet_beat~3 (
	.dataa(!\burst_uncompress_byte_counter[6]~q ),
	.datab(!\burst_uncompress_byte_counter[5]~q ),
	.datac(!\burst_uncompress_byte_counter[4]~q ),
	.datad(!\burst_uncompress_byte_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_packet_beat~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~3 .extended_lut = "off";
defparam \last_packet_beat~3 .lut_mask = 64'h8000800080008000;
defparam \last_packet_beat~3 .shared_arith = "off";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!mem_77_0),
	.datab(!mem_76_0),
	.datac(!mem_75_0),
	.datad(!mem_74_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h8000800080008000;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~6 (
	.dataa(!mem_78_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat2),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~6 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~6 .lut_mask = 64'h0000000C0A0A000C;
defparam \burst_uncompress_byte_counter~6 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[7] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[7]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[7] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[7] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[2]~q ),
	.datac(!\last_packet_beat~3_combout ),
	.datad(!\burst_uncompress_byte_counter[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~0 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~0 .lut_mask = 64'h5155515551555155;
defparam \burst_uncompress_byte_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!mem_77_0),
	.datab(!mem_76_0),
	.datac(!mem_75_0),
	.datad(!mem_74_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~2 (
	.dataa(!last_packet_beat2),
	.datab(!\burst_uncompress_byte_counter~0_combout ),
	.datac(!\Add0~1_combout ),
	.datad(!\Add1~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~2 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~2 .lut_mask = 64'h5410541054105410;
defparam \burst_uncompress_byte_counter~2 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[5] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[5]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[5] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[5] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h8000800080008000;
defparam \Add0~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~1 (
	.dataa(!mem_78_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat2),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~1 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~1 .lut_mask = 64'h0505030C0A0A030C;
defparam \burst_uncompress_byte_counter~1 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[6] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[6]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[6] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[6] .power_up = "low";

endmodule

module spw_babasu_altera_merlin_slave_agent_2 (
	waitrequest_reset_override,
	stateST_COMP_TRANS,
	out_valid_reg,
	mem_used_1,
	in_narrow_reg,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	WideOr0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	in_data_reg_68,
	cp_ready,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_129_0,
	mem_used_01,
	mem_66_0,
	comb,
	last_packet_beat,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	last_packet_beat1,
	altera_reset_synchronizer_int_chain_out,
	m0_write1,
	nxt_out_eop,
	cp_ready1,
	last_packet_beat2,
	WideOr01,
	read,
	cp_ready2,
	in_data_reg_69,
	rf_source_valid,
	rf_sink_ready,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	waitrequest_reset_override;
input 	stateST_COMP_TRANS;
input 	out_valid_reg;
input 	mem_used_1;
input 	in_narrow_reg;
input 	in_byteen_reg_3;
input 	in_byteen_reg_2;
input 	in_byteen_reg_1;
input 	in_byteen_reg_0;
output 	WideOr0;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	in_data_reg_68;
output 	cp_ready;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	mem_129_0;
input 	mem_used_01;
input 	mem_66_0;
output 	comb;
output 	last_packet_beat;
input 	mem_78_0;
input 	mem_77_0;
input 	mem_76_0;
input 	mem_75_0;
input 	mem_74_0;
output 	last_packet_beat1;
input 	altera_reset_synchronizer_int_chain_out;
output 	m0_write1;
input 	nxt_out_eop;
output 	cp_ready1;
output 	last_packet_beat2;
input 	WideOr01;
input 	read;
output 	cp_ready2;
input 	in_data_reg_69;
output 	rf_source_valid;
output 	rf_sink_ready;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \local_write~combout ;
wire \cp_ready~1_combout ;
wire \cp_ready~2_combout ;


spw_babasu_altera_merlin_burst_uncompressor_2 uncompressor(
	.mem_66_0(mem_66_0),
	.comb(comb),
	.last_packet_beat(last_packet_beat),
	.mem_78_0(mem_78_0),
	.mem_77_0(mem_77_0),
	.mem_76_0(mem_76_0),
	.mem_75_0(mem_75_0),
	.mem_74_0(mem_74_0),
	.last_packet_beat1(last_packet_beat1),
	.reset(altera_reset_synchronizer_int_chain_out),
	.last_packet_beat2(last_packet_beat2),
	.WideOr0(WideOr01),
	.read(read),
	.sink_ready(rf_sink_ready),
	.clk(clk_clk));

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!in_narrow_reg),
	.datac(!in_byteen_reg_3),
	.datad(!in_byteen_reg_2),
	.datae(!in_byteen_reg_1),
	.dataf(!in_byteen_reg_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h1FFFFFFFFFFFFFFF;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~0 (
	.dataa(!waitrequest_reset_override),
	.datab(!mem_used_1),
	.datac(!WideOr0),
	.datad(!wait_latency_counter_1),
	.datae(!wait_latency_counter_0),
	.dataf(!\local_write~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~0 .extended_lut = "off";
defparam \cp_ready~0 .lut_mask = 64'hC0C0C4C0C4C0C0C0;
defparam \cp_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \comb~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_129_0),
	.datad(!mem_used_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(comb),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~0 .extended_lut = "off";
defparam \comb~0 .lut_mask = 64'h007F007F007F007F;
defparam \comb~0 .shared_arith = "off";

cyclonev_lcell_comb m0_write(
	.dataa(!mem_used_1),
	.datab(!WideOr0),
	.datac(!\local_write~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write1),
	.sumout(),
	.cout(),
	.shareout());
defparam m0_write.extended_lut = "off";
defparam m0_write.lut_mask = 64'h0202020202020202;
defparam m0_write.shared_arith = "off";

cyclonev_lcell_comb \cp_ready~3 (
	.dataa(!mem_used_1),
	.datab(!in_narrow_reg),
	.datac(!\cp_ready~1_combout ),
	.datad(!\cp_ready~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~3 .extended_lut = "off";
defparam \cp_ready~3 .lut_mask = 64'h08AA08AA08AA08AA;
defparam \cp_ready~3 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~4 (
	.dataa(!waitrequest_reset_override),
	.datab(!mem_used_1),
	.datac(!WideOr0),
	.datad(!wait_latency_counter_1),
	.datae(!wait_latency_counter_0),
	.dataf(!\local_write~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready2),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~4 .extended_lut = "off";
defparam \cp_ready~4 .lut_mask = 64'h0000550004005100;
defparam \cp_ready~4 .shared_arith = "off";

cyclonev_lcell_comb \rf_source_valid~0 (
	.dataa(!in_data_reg_68),
	.datab(!out_valid_reg),
	.datac(!nxt_out_eop),
	.datad(!in_data_reg_69),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rf_source_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_source_valid~0 .extended_lut = "off";
defparam \rf_source_valid~0 .lut_mask = 64'h0133013301330133;
defparam \rf_source_valid~0 .shared_arith = "off";

cyclonev_lcell_comb local_write(
	.dataa(!in_data_reg_68),
	.datab(!out_valid_reg),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\local_write~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam local_write.extended_lut = "off";
defparam local_write.lut_mask = 64'h1111111111111111;
defparam local_write.shared_arith = "off";

cyclonev_lcell_comb \cp_ready~1 (
	.dataa(!in_byteen_reg_3),
	.datab(!in_byteen_reg_2),
	.datac(!in_byteen_reg_1),
	.datad(!in_byteen_reg_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cp_ready~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~1 .extended_lut = "off";
defparam \cp_ready~1 .lut_mask = 64'h8000800080008000;
defparam \cp_ready~1 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~2 (
	.dataa(!waitrequest_reset_override),
	.datab(!wait_latency_counter_1),
	.datac(!wait_latency_counter_0),
	.datad(!\local_write~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cp_ready~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~2 .extended_lut = "off";
defparam \cp_ready~2 .lut_mask = 64'h0440044004400440;
defparam \cp_ready~2 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_burst_uncompressor_2 (
	mem_66_0,
	comb,
	last_packet_beat,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	last_packet_beat1,
	reset,
	last_packet_beat2,
	WideOr0,
	read,
	sink_ready,
	clk)/* synthesis synthesis_greybox=0 */;
input 	mem_66_0;
input 	comb;
output 	last_packet_beat;
input 	mem_78_0;
input 	mem_77_0;
input 	mem_76_0;
input 	mem_75_0;
input 	mem_74_0;
output 	last_packet_beat1;
input 	reset;
output 	last_packet_beat2;
input 	WideOr0;
input 	read;
output 	sink_ready;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \burst_uncompress_busy~q ;
wire \burst_uncompress_byte_counter~5_combout ;
wire \burst_uncompress_byte_counter[2]~q ;
wire \burst_uncompress_byte_counter~4_combout ;
wire \burst_uncompress_byte_counter[3]~q ;
wire \Add0~2_combout ;
wire \burst_uncompress_byte_counter~3_combout ;
wire \burst_uncompress_byte_counter[4]~q ;
wire \last_packet_beat~3_combout ;
wire \Add1~0_combout ;
wire \burst_uncompress_byte_counter~6_combout ;
wire \burst_uncompress_byte_counter[7]~q ;
wire \burst_uncompress_byte_counter~0_combout ;
wire \Add0~1_combout ;
wire \Add1~1_combout ;
wire \burst_uncompress_byte_counter~2_combout ;
wire \burst_uncompress_byte_counter[5]~q ;
wire \Add0~0_combout ;
wire \burst_uncompress_byte_counter~1_combout ;
wire \burst_uncompress_byte_counter[6]~q ;


cyclonev_lcell_comb \last_packet_beat~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!\burst_uncompress_byte_counter[5]~q ),
	.datad(!\burst_uncompress_byte_counter[4]~q ),
	.datae(!\burst_uncompress_byte_counter[3]~q ),
	.dataf(!\burst_uncompress_byte_counter[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~0 .extended_lut = "off";
defparam \last_packet_beat~0 .lut_mask = 64'h0000000040000000;
defparam \last_packet_beat~0 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~1 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_78_0),
	.datac(!mem_77_0),
	.datad(!mem_76_0),
	.datae(!mem_75_0),
	.dataf(!mem_74_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat1),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~1 .extended_lut = "off";
defparam \last_packet_beat~1 .lut_mask = 64'h0000000080000000;
defparam \last_packet_beat~1 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~2 (
	.dataa(!comb),
	.datab(!mem_66_0),
	.datac(!last_packet_beat),
	.datad(!last_packet_beat1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat2),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~2 .extended_lut = "off";
defparam \last_packet_beat~2 .lut_mask = 64'h3222322232223222;
defparam \last_packet_beat~2 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!comb),
	.datad(!last_packet_beat2),
	.datae(!WideOr0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~0 .extended_lut = "off";
defparam \sink_ready~0 .lut_mask = 64'h00000F0000000F00;
defparam \sink_ready~0 .shared_arith = "off";

dffeas burst_uncompress_busy(
	.clk(clk),
	.d(last_packet_beat2),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_busy~q ),
	.prn(vcc));
defparam burst_uncompress_busy.is_wysiwyg = "true";
defparam burst_uncompress_busy.power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~5 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_74_0),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(!last_packet_beat2),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~5 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~5 .lut_mask = 64'h00C800FA00C800FA;
defparam \burst_uncompress_byte_counter~5 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[2] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[2]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[2] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[2] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~4 (
	.dataa(!mem_75_0),
	.datab(!mem_74_0),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(!last_packet_beat2),
	.dataf(!\burst_uncompress_byte_counter~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~4 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~4 .lut_mask = 64'h000099990000F00F;
defparam \burst_uncompress_byte_counter~4 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[3] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[3]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[3] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[3] .power_up = "low";

cyclonev_lcell_comb \Add0~2 (
	.dataa(!\burst_uncompress_byte_counter[4]~q ),
	.datab(!\burst_uncompress_byte_counter[3]~q ),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~2 .extended_lut = "off";
defparam \Add0~2 .lut_mask = 64'h6A6A6A6A6A6A6A6A;
defparam \Add0~2 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~3 (
	.dataa(!mem_76_0),
	.datab(!mem_75_0),
	.datac(!mem_74_0),
	.datad(!last_packet_beat2),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add0~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~3 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~3 .lut_mask = 64'h009500FF00950000;
defparam \burst_uncompress_byte_counter~3 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[4] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[4]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[4] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[4] .power_up = "low";

cyclonev_lcell_comb \last_packet_beat~3 (
	.dataa(!\burst_uncompress_byte_counter[6]~q ),
	.datab(!\burst_uncompress_byte_counter[5]~q ),
	.datac(!\burst_uncompress_byte_counter[4]~q ),
	.datad(!\burst_uncompress_byte_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_packet_beat~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~3 .extended_lut = "off";
defparam \last_packet_beat~3 .lut_mask = 64'h8000800080008000;
defparam \last_packet_beat~3 .shared_arith = "off";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!mem_77_0),
	.datab(!mem_76_0),
	.datac(!mem_75_0),
	.datad(!mem_74_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h8000800080008000;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~6 (
	.dataa(!mem_78_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat2),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~6 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~6 .lut_mask = 64'h0000000C0A0A000C;
defparam \burst_uncompress_byte_counter~6 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[7] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[7]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[7] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[7] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[2]~q ),
	.datac(!\last_packet_beat~3_combout ),
	.datad(!\burst_uncompress_byte_counter[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~0 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~0 .lut_mask = 64'h5155515551555155;
defparam \burst_uncompress_byte_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!mem_77_0),
	.datab(!mem_76_0),
	.datac(!mem_75_0),
	.datad(!mem_74_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~2 (
	.dataa(!last_packet_beat2),
	.datab(!\burst_uncompress_byte_counter~0_combout ),
	.datac(!\Add0~1_combout ),
	.datad(!\Add1~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~2 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~2 .lut_mask = 64'h5410541054105410;
defparam \burst_uncompress_byte_counter~2 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[5] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[5]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[5] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[5] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h8000800080008000;
defparam \Add0~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~1 (
	.dataa(!mem_78_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat2),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~1 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~1 .lut_mask = 64'h0505030C0A0A030C;
defparam \burst_uncompress_byte_counter~1 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[6] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[6]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[6] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[6] .power_up = "low";

endmodule

module spw_babasu_altera_merlin_slave_agent_3 (
	h2f_RREADY_0,
	stateST_COMP_TRANS,
	mem_used_1,
	waitrequest_reset_override,
	in_data_reg_69,
	in_narrow_reg,
	wait_latency_counter_1,
	wait_latency_counter_0,
	cp_ready,
	cp_ready1,
	empty,
	mem_66_0,
	mem_used_0,
	last_packet_beat,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	last_packet_beat1,
	altera_reset_synchronizer_int_chain_out,
	last_packet_beat2,
	cp_ready2,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_RREADY_0;
input 	stateST_COMP_TRANS;
input 	mem_used_1;
input 	waitrequest_reset_override;
input 	in_data_reg_69;
input 	in_narrow_reg;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
output 	cp_ready;
output 	cp_ready1;
input 	empty;
input 	mem_66_0;
input 	mem_used_0;
output 	last_packet_beat;
input 	mem_78_0;
input 	mem_77_0;
input 	mem_76_0;
input 	mem_75_0;
input 	mem_74_0;
output 	last_packet_beat1;
input 	altera_reset_synchronizer_int_chain_out;
output 	last_packet_beat2;
output 	cp_ready2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



spw_babasu_altera_merlin_burst_uncompressor_3 uncompressor(
	.h2f_RREADY_0(h2f_RREADY_0),
	.empty(empty),
	.mem_66_0(mem_66_0),
	.mem_used_0(mem_used_0),
	.last_packet_beat(last_packet_beat),
	.mem_78_0(mem_78_0),
	.mem_77_0(mem_77_0),
	.mem_76_0(mem_76_0),
	.mem_75_0(mem_75_0),
	.mem_74_0(mem_74_0),
	.last_packet_beat1(last_packet_beat1),
	.reset(altera_reset_synchronizer_int_chain_out),
	.last_packet_beat2(last_packet_beat2),
	.clk(clk_clk));

cyclonev_lcell_comb \cp_ready~0 (
	.dataa(!waitrequest_reset_override),
	.datab(!in_data_reg_69),
	.datac(!stateST_COMP_TRANS),
	.datad(!in_narrow_reg),
	.datae(!wait_latency_counter_1),
	.dataf(!wait_latency_counter_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~0 .extended_lut = "off";
defparam \cp_ready~0 .lut_mask = 64'hCCC0CCC0DDD5CCC0;
defparam \cp_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~1 (
	.dataa(!mem_used_1),
	.datab(!cp_ready),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~1 .extended_lut = "off";
defparam \cp_ready~1 .lut_mask = 64'h2222222222222222;
defparam \cp_ready~1 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~2 (
	.dataa(!waitrequest_reset_override),
	.datab(!in_data_reg_69),
	.datac(!in_narrow_reg),
	.datad(!wait_latency_counter_1),
	.datae(!wait_latency_counter_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready2),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~2 .extended_lut = "off";
defparam \cp_ready~2 .lut_mask = 64'hC0C0D5C0C0C0D5C0;
defparam \cp_ready~2 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_burst_uncompressor_3 (
	h2f_RREADY_0,
	empty,
	mem_66_0,
	mem_used_0,
	last_packet_beat,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	last_packet_beat1,
	reset,
	last_packet_beat2,
	clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_RREADY_0;
input 	empty;
input 	mem_66_0;
input 	mem_used_0;
output 	last_packet_beat;
input 	mem_78_0;
input 	mem_77_0;
input 	mem_76_0;
input 	mem_75_0;
input 	mem_74_0;
output 	last_packet_beat1;
input 	reset;
output 	last_packet_beat2;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always0~0_combout ;
wire \burst_uncompress_busy~q ;
wire \burst_uncompress_byte_counter~5_combout ;
wire \burst_uncompress_byte_counter[2]~q ;
wire \burst_uncompress_byte_counter~4_combout ;
wire \burst_uncompress_byte_counter[3]~q ;
wire \Add0~2_combout ;
wire \burst_uncompress_byte_counter~3_combout ;
wire \burst_uncompress_byte_counter[4]~q ;
wire \last_packet_beat~3_combout ;
wire \Add1~0_combout ;
wire \burst_uncompress_byte_counter~6_combout ;
wire \burst_uncompress_byte_counter[7]~q ;
wire \burst_uncompress_byte_counter~0_combout ;
wire \Add0~1_combout ;
wire \Add1~1_combout ;
wire \burst_uncompress_byte_counter~2_combout ;
wire \burst_uncompress_byte_counter[5]~q ;
wire \Add0~0_combout ;
wire \burst_uncompress_byte_counter~1_combout ;
wire \burst_uncompress_byte_counter[6]~q ;


cyclonev_lcell_comb \last_packet_beat~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!\burst_uncompress_byte_counter[5]~q ),
	.datad(!\burst_uncompress_byte_counter[4]~q ),
	.datae(!\burst_uncompress_byte_counter[3]~q ),
	.dataf(!\burst_uncompress_byte_counter[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~0 .extended_lut = "off";
defparam \last_packet_beat~0 .lut_mask = 64'h0000000040000000;
defparam \last_packet_beat~0 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~1 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_78_0),
	.datac(!mem_77_0),
	.datad(!mem_76_0),
	.datae(!mem_75_0),
	.dataf(!mem_74_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat1),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~1 .extended_lut = "off";
defparam \last_packet_beat~1 .lut_mask = 64'h0000000080000000;
defparam \last_packet_beat~1 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~2 (
	.dataa(!empty),
	.datab(!mem_66_0),
	.datac(!mem_used_0),
	.datad(!last_packet_beat),
	.datae(!last_packet_beat1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat2),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~2 .extended_lut = "off";
defparam \last_packet_beat~2 .lut_mask = 64'h3331313133313131;
defparam \last_packet_beat~2 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!h2f_RREADY_0),
	.datab(!empty),
	.datac(!mem_used_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'h0404040404040404;
defparam \always0~0 .shared_arith = "off";

dffeas burst_uncompress_busy(
	.clk(clk),
	.d(last_packet_beat2),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_busy~q ),
	.prn(vcc));
defparam burst_uncompress_busy.is_wysiwyg = "true";
defparam burst_uncompress_busy.power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~5 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_74_0),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(!last_packet_beat2),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~5 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~5 .lut_mask = 64'h00C800FA00C800FA;
defparam \burst_uncompress_byte_counter~5 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[2] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[2]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[2] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[2] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~4 (
	.dataa(!mem_75_0),
	.datab(!mem_74_0),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(!last_packet_beat2),
	.dataf(!\burst_uncompress_byte_counter~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~4 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~4 .lut_mask = 64'h000099990000F00F;
defparam \burst_uncompress_byte_counter~4 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[3] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[3]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[3] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[3] .power_up = "low";

cyclonev_lcell_comb \Add0~2 (
	.dataa(!\burst_uncompress_byte_counter[4]~q ),
	.datab(!\burst_uncompress_byte_counter[3]~q ),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~2 .extended_lut = "off";
defparam \Add0~2 .lut_mask = 64'h6A6A6A6A6A6A6A6A;
defparam \Add0~2 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~3 (
	.dataa(!mem_76_0),
	.datab(!mem_75_0),
	.datac(!mem_74_0),
	.datad(!last_packet_beat2),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add0~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~3 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~3 .lut_mask = 64'h009500FF00950000;
defparam \burst_uncompress_byte_counter~3 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[4] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[4]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[4] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[4] .power_up = "low";

cyclonev_lcell_comb \last_packet_beat~3 (
	.dataa(!\burst_uncompress_byte_counter[6]~q ),
	.datab(!\burst_uncompress_byte_counter[5]~q ),
	.datac(!\burst_uncompress_byte_counter[4]~q ),
	.datad(!\burst_uncompress_byte_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_packet_beat~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~3 .extended_lut = "off";
defparam \last_packet_beat~3 .lut_mask = 64'h8000800080008000;
defparam \last_packet_beat~3 .shared_arith = "off";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!mem_77_0),
	.datab(!mem_76_0),
	.datac(!mem_75_0),
	.datad(!mem_74_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h8000800080008000;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~6 (
	.dataa(!mem_78_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat2),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~6 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~6 .lut_mask = 64'h0000000C0A0A000C;
defparam \burst_uncompress_byte_counter~6 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[7] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[7]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[7] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[7] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[2]~q ),
	.datac(!\last_packet_beat~3_combout ),
	.datad(!\burst_uncompress_byte_counter[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~0 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~0 .lut_mask = 64'h5155515551555155;
defparam \burst_uncompress_byte_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!mem_77_0),
	.datab(!mem_76_0),
	.datac(!mem_75_0),
	.datad(!mem_74_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~2 (
	.dataa(!last_packet_beat2),
	.datab(!\burst_uncompress_byte_counter~0_combout ),
	.datac(!\Add0~1_combout ),
	.datad(!\Add1~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~2 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~2 .lut_mask = 64'h5410541054105410;
defparam \burst_uncompress_byte_counter~2 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[5] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[5]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[5] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[5] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h8000800080008000;
defparam \Add0~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~1 (
	.dataa(!mem_78_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat2),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~1 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~1 .lut_mask = 64'h0505030C0A0A030C;
defparam \burst_uncompress_byte_counter~1 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[6] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[6]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[6] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[6] .power_up = "low";

endmodule

module spw_babasu_altera_merlin_slave_agent_4 (
	h2f_RREADY_0,
	waitrequest_reset_override,
	in_data_reg_69,
	stateST_COMP_TRANS,
	in_narrow_reg,
	wait_latency_counter_1,
	wait_latency_counter_0,
	cp_ready,
	empty,
	mem_66_0,
	mem_used_0,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	last_packet_beat,
	altera_reset_synchronizer_int_chain_out,
	cp_ready1,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_RREADY_0;
input 	waitrequest_reset_override;
input 	in_data_reg_69;
input 	stateST_COMP_TRANS;
input 	in_narrow_reg;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
output 	cp_ready;
input 	empty;
input 	mem_66_0;
input 	mem_used_0;
input 	mem_78_0;
input 	mem_77_0;
input 	mem_76_0;
input 	mem_75_0;
input 	mem_74_0;
output 	last_packet_beat;
input 	altera_reset_synchronizer_int_chain_out;
output 	cp_ready1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



spw_babasu_altera_merlin_burst_uncompressor_4 uncompressor(
	.h2f_RREADY_0(h2f_RREADY_0),
	.empty(empty),
	.mem_66_0(mem_66_0),
	.mem_used_0(mem_used_0),
	.mem_78_0(mem_78_0),
	.mem_77_0(mem_77_0),
	.mem_76_0(mem_76_0),
	.mem_75_0(mem_75_0),
	.mem_74_0(mem_74_0),
	.last_packet_beat(last_packet_beat),
	.reset(altera_reset_synchronizer_int_chain_out),
	.clk(clk_clk));

cyclonev_lcell_comb \cp_ready~0 (
	.dataa(!waitrequest_reset_override),
	.datab(!in_data_reg_69),
	.datac(!stateST_COMP_TRANS),
	.datad(!in_narrow_reg),
	.datae(!wait_latency_counter_1),
	.dataf(!wait_latency_counter_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~0 .extended_lut = "off";
defparam \cp_ready~0 .lut_mask = 64'hCCC0CCC0DDD5CCC0;
defparam \cp_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~1 (
	.dataa(!waitrequest_reset_override),
	.datab(!in_data_reg_69),
	.datac(!in_narrow_reg),
	.datad(!wait_latency_counter_1),
	.datae(!wait_latency_counter_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~1 .extended_lut = "off";
defparam \cp_ready~1 .lut_mask = 64'hC0C0D5C0C0C0D5C0;
defparam \cp_ready~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_burst_uncompressor_4 (
	h2f_RREADY_0,
	empty,
	mem_66_0,
	mem_used_0,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	last_packet_beat,
	reset,
	clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_RREADY_0;
input 	empty;
input 	mem_66_0;
input 	mem_used_0;
input 	mem_78_0;
input 	mem_77_0;
input 	mem_76_0;
input 	mem_75_0;
input 	mem_74_0;
output 	last_packet_beat;
input 	reset;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always0~0_combout ;
wire \burst_uncompress_busy~q ;
wire \burst_uncompress_byte_counter~5_combout ;
wire \burst_uncompress_byte_counter[3]~q ;
wire \Add0~2_combout ;
wire \burst_uncompress_byte_counter~4_combout ;
wire \burst_uncompress_byte_counter[4]~q ;
wire \Add0~1_combout ;
wire \Add1~1_combout ;
wire \burst_uncompress_byte_counter~3_combout ;
wire \burst_uncompress_byte_counter[5]~q ;
wire \Add0~0_combout ;
wire \Add1~0_combout ;
wire \burst_uncompress_byte_counter~2_combout ;
wire \burst_uncompress_byte_counter[6]~q ;
wire \last_packet_beat~1_combout ;
wire \burst_uncompress_byte_counter~6_combout ;
wire \burst_uncompress_byte_counter[7]~q ;
wire \burst_uncompress_byte_counter~0_combout ;
wire \burst_uncompress_byte_counter~1_combout ;
wire \burst_uncompress_byte_counter[2]~q ;
wire \last_packet_beat~0_combout ;
wire \last_packet_beat~2_combout ;


cyclonev_lcell_comb \last_packet_beat~3 (
	.dataa(!empty),
	.datab(!mem_66_0),
	.datac(!mem_used_0),
	.datad(!\last_packet_beat~0_combout ),
	.datae(!\last_packet_beat~1_combout ),
	.dataf(!\last_packet_beat~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~3 .extended_lut = "off";
defparam \last_packet_beat~3 .lut_mask = 64'h3333333131313131;
defparam \last_packet_beat~3 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!h2f_RREADY_0),
	.datab(!empty),
	.datac(!mem_used_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'h0404040404040404;
defparam \always0~0 .shared_arith = "off";

dffeas burst_uncompress_busy(
	.clk(clk),
	.d(last_packet_beat),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_busy~q ),
	.prn(vcc));
defparam burst_uncompress_busy.is_wysiwyg = "true";
defparam burst_uncompress_busy.power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~5 (
	.dataa(!mem_75_0),
	.datab(!mem_74_0),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(!last_packet_beat),
	.dataf(!\burst_uncompress_byte_counter~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~5 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~5 .lut_mask = 64'h000099990000F00F;
defparam \burst_uncompress_byte_counter~5 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[3] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[3]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[3] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[3] .power_up = "low";

cyclonev_lcell_comb \Add0~2 (
	.dataa(!\burst_uncompress_byte_counter[4]~q ),
	.datab(!\burst_uncompress_byte_counter[3]~q ),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~2 .extended_lut = "off";
defparam \Add0~2 .lut_mask = 64'h6A6A6A6A6A6A6A6A;
defparam \Add0~2 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~4 (
	.dataa(!mem_76_0),
	.datab(!mem_75_0),
	.datac(!mem_74_0),
	.datad(!last_packet_beat),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add0~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~4 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~4 .lut_mask = 64'h009500FF00950000;
defparam \burst_uncompress_byte_counter~4 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[4] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[4]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[4] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[4] .power_up = "low";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!mem_77_0),
	.datab(!mem_76_0),
	.datac(!mem_75_0),
	.datad(!mem_74_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~3 (
	.dataa(!last_packet_beat),
	.datab(!\burst_uncompress_byte_counter~0_combout ),
	.datac(!\Add0~1_combout ),
	.datad(!\Add1~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~3 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~3 .lut_mask = 64'h5410541054105410;
defparam \burst_uncompress_byte_counter~3 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[5] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[5]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[5] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[5] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h8000800080008000;
defparam \Add0~0 .shared_arith = "off";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!mem_77_0),
	.datab(!mem_76_0),
	.datac(!mem_75_0),
	.datad(!mem_74_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h8000800080008000;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~2 (
	.dataa(!mem_78_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~2 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~2 .lut_mask = 64'h0505030C0A0A030C;
defparam \burst_uncompress_byte_counter~2 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[6] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[6]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[6] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[6] .power_up = "low";

cyclonev_lcell_comb \last_packet_beat~1 (
	.dataa(!\burst_uncompress_byte_counter[6]~q ),
	.datab(!\burst_uncompress_byte_counter[5]~q ),
	.datac(!\burst_uncompress_byte_counter[4]~q ),
	.datad(!\burst_uncompress_byte_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_packet_beat~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~1 .extended_lut = "off";
defparam \last_packet_beat~1 .lut_mask = 64'h8000800080008000;
defparam \last_packet_beat~1 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~6 (
	.dataa(!mem_78_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~6 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~6 .lut_mask = 64'h0000000C0A0A000C;
defparam \burst_uncompress_byte_counter~6 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[7] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[7]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[7] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[7] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[2]~q ),
	.datac(!\last_packet_beat~1_combout ),
	.datad(!\burst_uncompress_byte_counter[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~0 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~0 .lut_mask = 64'h5155515551555155;
defparam \burst_uncompress_byte_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~1 (
	.dataa(!mem_74_0),
	.datab(!\last_packet_beat~0_combout ),
	.datac(!last_packet_beat),
	.datad(!\burst_uncompress_byte_counter~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~1 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~1 .lut_mask = 64'h080C080C080C080C;
defparam \burst_uncompress_byte_counter~1 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[2] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[2]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[2] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[2] .power_up = "low";

cyclonev_lcell_comb \last_packet_beat~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_packet_beat~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~0 .extended_lut = "off";
defparam \last_packet_beat~0 .lut_mask = 64'h1111111111111111;
defparam \last_packet_beat~0 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~2 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_78_0),
	.datac(!mem_77_0),
	.datad(!mem_76_0),
	.datae(!mem_75_0),
	.dataf(!mem_74_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_packet_beat~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~2 .extended_lut = "off";
defparam \last_packet_beat~2 .lut_mask = 64'h0000000080000000;
defparam \last_packet_beat~2 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_slave_agent_5 (
	waitrequest_reset_override,
	stateST_COMP_TRANS,
	out_valid_reg,
	mem_used_1,
	in_narrow_reg,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	WideOr0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	in_data_reg_68,
	cp_ready,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_129_0,
	mem_used_01,
	mem_66_0,
	comb,
	last_packet_beat,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	last_packet_beat1,
	altera_reset_synchronizer_int_chain_out,
	m0_write1,
	nxt_out_eop,
	cp_ready1,
	last_packet_beat2,
	WideOr01,
	read,
	cp_ready2,
	in_data_reg_69,
	rf_source_valid,
	rf_sink_ready,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	waitrequest_reset_override;
input 	stateST_COMP_TRANS;
input 	out_valid_reg;
input 	mem_used_1;
input 	in_narrow_reg;
input 	in_byteen_reg_3;
input 	in_byteen_reg_2;
input 	in_byteen_reg_1;
input 	in_byteen_reg_0;
output 	WideOr0;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	in_data_reg_68;
output 	cp_ready;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	mem_129_0;
input 	mem_used_01;
input 	mem_66_0;
output 	comb;
output 	last_packet_beat;
input 	mem_78_0;
input 	mem_77_0;
input 	mem_76_0;
input 	mem_75_0;
input 	mem_74_0;
output 	last_packet_beat1;
input 	altera_reset_synchronizer_int_chain_out;
output 	m0_write1;
input 	nxt_out_eop;
output 	cp_ready1;
output 	last_packet_beat2;
input 	WideOr01;
input 	read;
output 	cp_ready2;
input 	in_data_reg_69;
output 	rf_source_valid;
output 	rf_sink_ready;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \local_write~combout ;
wire \cp_ready~1_combout ;
wire \cp_ready~2_combout ;


spw_babasu_altera_merlin_burst_uncompressor_5 uncompressor(
	.mem_66_0(mem_66_0),
	.comb(comb),
	.last_packet_beat(last_packet_beat),
	.mem_78_0(mem_78_0),
	.mem_77_0(mem_77_0),
	.mem_76_0(mem_76_0),
	.mem_75_0(mem_75_0),
	.mem_74_0(mem_74_0),
	.last_packet_beat1(last_packet_beat1),
	.reset(altera_reset_synchronizer_int_chain_out),
	.last_packet_beat2(last_packet_beat2),
	.WideOr0(WideOr01),
	.read(read),
	.sink_ready(rf_sink_ready),
	.clk(clk_clk));

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!in_narrow_reg),
	.datac(!in_byteen_reg_3),
	.datad(!in_byteen_reg_2),
	.datae(!in_byteen_reg_1),
	.dataf(!in_byteen_reg_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h1FFFFFFFFFFFFFFF;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~0 (
	.dataa(!waitrequest_reset_override),
	.datab(!mem_used_1),
	.datac(!WideOr0),
	.datad(!wait_latency_counter_1),
	.datae(!wait_latency_counter_0),
	.dataf(!\local_write~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~0 .extended_lut = "off";
defparam \cp_ready~0 .lut_mask = 64'hC0C0C4C0C4C0C0C0;
defparam \cp_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \comb~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_129_0),
	.datad(!mem_used_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(comb),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~0 .extended_lut = "off";
defparam \comb~0 .lut_mask = 64'h007F007F007F007F;
defparam \comb~0 .shared_arith = "off";

cyclonev_lcell_comb m0_write(
	.dataa(!mem_used_1),
	.datab(!WideOr0),
	.datac(!\local_write~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write1),
	.sumout(),
	.cout(),
	.shareout());
defparam m0_write.extended_lut = "off";
defparam m0_write.lut_mask = 64'h0202020202020202;
defparam m0_write.shared_arith = "off";

cyclonev_lcell_comb \cp_ready~3 (
	.dataa(!mem_used_1),
	.datab(!in_narrow_reg),
	.datac(!\cp_ready~1_combout ),
	.datad(!\cp_ready~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~3 .extended_lut = "off";
defparam \cp_ready~3 .lut_mask = 64'h08AA08AA08AA08AA;
defparam \cp_ready~3 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~4 (
	.dataa(!waitrequest_reset_override),
	.datab(!mem_used_1),
	.datac(!WideOr0),
	.datad(!wait_latency_counter_1),
	.datae(!wait_latency_counter_0),
	.dataf(!\local_write~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready2),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~4 .extended_lut = "off";
defparam \cp_ready~4 .lut_mask = 64'h0000550004005100;
defparam \cp_ready~4 .shared_arith = "off";

cyclonev_lcell_comb \rf_source_valid~0 (
	.dataa(!in_data_reg_68),
	.datab(!out_valid_reg),
	.datac(!nxt_out_eop),
	.datad(!in_data_reg_69),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rf_source_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_source_valid~0 .extended_lut = "off";
defparam \rf_source_valid~0 .lut_mask = 64'h0133013301330133;
defparam \rf_source_valid~0 .shared_arith = "off";

cyclonev_lcell_comb local_write(
	.dataa(!in_data_reg_68),
	.datab(!out_valid_reg),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\local_write~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam local_write.extended_lut = "off";
defparam local_write.lut_mask = 64'h1111111111111111;
defparam local_write.shared_arith = "off";

cyclonev_lcell_comb \cp_ready~1 (
	.dataa(!in_byteen_reg_3),
	.datab(!in_byteen_reg_2),
	.datac(!in_byteen_reg_1),
	.datad(!in_byteen_reg_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cp_ready~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~1 .extended_lut = "off";
defparam \cp_ready~1 .lut_mask = 64'h8000800080008000;
defparam \cp_ready~1 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~2 (
	.dataa(!waitrequest_reset_override),
	.datab(!wait_latency_counter_1),
	.datac(!wait_latency_counter_0),
	.datad(!\local_write~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cp_ready~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~2 .extended_lut = "off";
defparam \cp_ready~2 .lut_mask = 64'h0440044004400440;
defparam \cp_ready~2 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_burst_uncompressor_5 (
	mem_66_0,
	comb,
	last_packet_beat,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	last_packet_beat1,
	reset,
	last_packet_beat2,
	WideOr0,
	read,
	sink_ready,
	clk)/* synthesis synthesis_greybox=0 */;
input 	mem_66_0;
input 	comb;
output 	last_packet_beat;
input 	mem_78_0;
input 	mem_77_0;
input 	mem_76_0;
input 	mem_75_0;
input 	mem_74_0;
output 	last_packet_beat1;
input 	reset;
output 	last_packet_beat2;
input 	WideOr0;
input 	read;
output 	sink_ready;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \burst_uncompress_busy~q ;
wire \burst_uncompress_byte_counter~5_combout ;
wire \burst_uncompress_byte_counter[2]~q ;
wire \burst_uncompress_byte_counter~4_combout ;
wire \burst_uncompress_byte_counter[3]~q ;
wire \Add0~2_combout ;
wire \burst_uncompress_byte_counter~3_combout ;
wire \burst_uncompress_byte_counter[4]~q ;
wire \last_packet_beat~3_combout ;
wire \Add1~0_combout ;
wire \burst_uncompress_byte_counter~6_combout ;
wire \burst_uncompress_byte_counter[7]~q ;
wire \burst_uncompress_byte_counter~0_combout ;
wire \Add0~1_combout ;
wire \Add1~1_combout ;
wire \burst_uncompress_byte_counter~2_combout ;
wire \burst_uncompress_byte_counter[5]~q ;
wire \Add0~0_combout ;
wire \burst_uncompress_byte_counter~1_combout ;
wire \burst_uncompress_byte_counter[6]~q ;


cyclonev_lcell_comb \last_packet_beat~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!\burst_uncompress_byte_counter[5]~q ),
	.datad(!\burst_uncompress_byte_counter[4]~q ),
	.datae(!\burst_uncompress_byte_counter[3]~q ),
	.dataf(!\burst_uncompress_byte_counter[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~0 .extended_lut = "off";
defparam \last_packet_beat~0 .lut_mask = 64'h0000000040000000;
defparam \last_packet_beat~0 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~1 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_78_0),
	.datac(!mem_77_0),
	.datad(!mem_76_0),
	.datae(!mem_75_0),
	.dataf(!mem_74_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat1),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~1 .extended_lut = "off";
defparam \last_packet_beat~1 .lut_mask = 64'h0000000080000000;
defparam \last_packet_beat~1 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~2 (
	.dataa(!comb),
	.datab(!mem_66_0),
	.datac(!last_packet_beat),
	.datad(!last_packet_beat1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat2),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~2 .extended_lut = "off";
defparam \last_packet_beat~2 .lut_mask = 64'h3222322232223222;
defparam \last_packet_beat~2 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!comb),
	.datad(!last_packet_beat2),
	.datae(!WideOr0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~0 .extended_lut = "off";
defparam \sink_ready~0 .lut_mask = 64'h00000F0000000F00;
defparam \sink_ready~0 .shared_arith = "off";

dffeas burst_uncompress_busy(
	.clk(clk),
	.d(last_packet_beat2),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_busy~q ),
	.prn(vcc));
defparam burst_uncompress_busy.is_wysiwyg = "true";
defparam burst_uncompress_busy.power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~5 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_74_0),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(!last_packet_beat2),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~5 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~5 .lut_mask = 64'h00C800FA00C800FA;
defparam \burst_uncompress_byte_counter~5 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[2] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[2]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[2] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[2] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~4 (
	.dataa(!mem_75_0),
	.datab(!mem_74_0),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(!last_packet_beat2),
	.dataf(!\burst_uncompress_byte_counter~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~4 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~4 .lut_mask = 64'h000099990000F00F;
defparam \burst_uncompress_byte_counter~4 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[3] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[3]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[3] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[3] .power_up = "low";

cyclonev_lcell_comb \Add0~2 (
	.dataa(!\burst_uncompress_byte_counter[4]~q ),
	.datab(!\burst_uncompress_byte_counter[3]~q ),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~2 .extended_lut = "off";
defparam \Add0~2 .lut_mask = 64'h6A6A6A6A6A6A6A6A;
defparam \Add0~2 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~3 (
	.dataa(!mem_76_0),
	.datab(!mem_75_0),
	.datac(!mem_74_0),
	.datad(!last_packet_beat2),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add0~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~3 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~3 .lut_mask = 64'h009500FF00950000;
defparam \burst_uncompress_byte_counter~3 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[4] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[4]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[4] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[4] .power_up = "low";

cyclonev_lcell_comb \last_packet_beat~3 (
	.dataa(!\burst_uncompress_byte_counter[6]~q ),
	.datab(!\burst_uncompress_byte_counter[5]~q ),
	.datac(!\burst_uncompress_byte_counter[4]~q ),
	.datad(!\burst_uncompress_byte_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_packet_beat~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~3 .extended_lut = "off";
defparam \last_packet_beat~3 .lut_mask = 64'h8000800080008000;
defparam \last_packet_beat~3 .shared_arith = "off";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!mem_77_0),
	.datab(!mem_76_0),
	.datac(!mem_75_0),
	.datad(!mem_74_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h8000800080008000;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~6 (
	.dataa(!mem_78_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat2),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~6 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~6 .lut_mask = 64'h0000000C0A0A000C;
defparam \burst_uncompress_byte_counter~6 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[7] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[7]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[7] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[7] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[2]~q ),
	.datac(!\last_packet_beat~3_combout ),
	.datad(!\burst_uncompress_byte_counter[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~0 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~0 .lut_mask = 64'h5155515551555155;
defparam \burst_uncompress_byte_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!mem_77_0),
	.datab(!mem_76_0),
	.datac(!mem_75_0),
	.datad(!mem_74_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~2 (
	.dataa(!last_packet_beat2),
	.datab(!\burst_uncompress_byte_counter~0_combout ),
	.datac(!\Add0~1_combout ),
	.datad(!\Add1~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~2 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~2 .lut_mask = 64'h5410541054105410;
defparam \burst_uncompress_byte_counter~2 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[5] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[5]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[5] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[5] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h8000800080008000;
defparam \Add0~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~1 (
	.dataa(!mem_78_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat2),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~1 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~1 .lut_mask = 64'h0505030C0A0A030C;
defparam \burst_uncompress_byte_counter~1 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[6] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[6]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[6] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[6] .power_up = "low";

endmodule

module spw_babasu_altera_merlin_slave_agent_6 (
	waitrequest_reset_override,
	stateST_COMP_TRANS,
	out_valid_reg,
	mem_used_1,
	in_narrow_reg,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	WideOr0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	in_data_reg_68,
	cp_ready,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_129_0,
	mem_used_01,
	mem_66_0,
	comb,
	last_packet_beat,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	last_packet_beat1,
	altera_reset_synchronizer_int_chain_out,
	m0_write1,
	nxt_out_eop,
	cp_ready1,
	last_packet_beat2,
	WideOr01,
	read,
	cp_ready2,
	in_data_reg_69,
	rf_source_valid,
	rf_sink_ready,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	waitrequest_reset_override;
input 	stateST_COMP_TRANS;
input 	out_valid_reg;
input 	mem_used_1;
input 	in_narrow_reg;
input 	in_byteen_reg_3;
input 	in_byteen_reg_2;
input 	in_byteen_reg_1;
input 	in_byteen_reg_0;
output 	WideOr0;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	in_data_reg_68;
output 	cp_ready;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	mem_129_0;
input 	mem_used_01;
input 	mem_66_0;
output 	comb;
output 	last_packet_beat;
input 	mem_78_0;
input 	mem_77_0;
input 	mem_76_0;
input 	mem_75_0;
input 	mem_74_0;
output 	last_packet_beat1;
input 	altera_reset_synchronizer_int_chain_out;
output 	m0_write1;
input 	nxt_out_eop;
output 	cp_ready1;
output 	last_packet_beat2;
input 	WideOr01;
input 	read;
output 	cp_ready2;
input 	in_data_reg_69;
output 	rf_source_valid;
output 	rf_sink_ready;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \local_write~combout ;
wire \cp_ready~1_combout ;


spw_babasu_altera_merlin_burst_uncompressor_6 uncompressor(
	.mem_66_0(mem_66_0),
	.comb(comb),
	.last_packet_beat(last_packet_beat),
	.mem_78_0(mem_78_0),
	.mem_77_0(mem_77_0),
	.mem_76_0(mem_76_0),
	.mem_75_0(mem_75_0),
	.mem_74_0(mem_74_0),
	.last_packet_beat1(last_packet_beat1),
	.reset(altera_reset_synchronizer_int_chain_out),
	.last_packet_beat2(last_packet_beat2),
	.WideOr0(WideOr01),
	.read(read),
	.sink_ready(rf_sink_ready),
	.clk(clk_clk));

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!in_narrow_reg),
	.datac(!in_byteen_reg_3),
	.datad(!in_byteen_reg_2),
	.datae(!in_byteen_reg_1),
	.dataf(!in_byteen_reg_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h1FFFFFFFFFFFFFFF;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~0 (
	.dataa(!mem_used_1),
	.datab(!WideOr0),
	.datac(!waitrequest_reset_override),
	.datad(!wait_latency_counter_1),
	.datae(!wait_latency_counter_0),
	.dataf(!\local_write~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~0 .extended_lut = "off";
defparam \cp_ready~0 .lut_mask = 64'h88888A888A888888;
defparam \cp_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \comb~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_129_0),
	.datad(!mem_used_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(comb),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~0 .extended_lut = "off";
defparam \comb~0 .lut_mask = 64'h007F007F007F007F;
defparam \comb~0 .shared_arith = "off";

cyclonev_lcell_comb m0_write(
	.dataa(!mem_used_1),
	.datab(!WideOr0),
	.datac(!\local_write~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write1),
	.sumout(),
	.cout(),
	.shareout());
defparam m0_write.extended_lut = "off";
defparam m0_write.lut_mask = 64'h0202020202020202;
defparam m0_write.shared_arith = "off";

cyclonev_lcell_comb \cp_ready~2 (
	.dataa(!waitrequest_reset_override),
	.datab(!wait_latency_counter_1),
	.datac(!wait_latency_counter_0),
	.datad(!\local_write~combout ),
	.datae(!\cp_ready~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~2 .extended_lut = "off";
defparam \cp_ready~2 .lut_mask = 64'hFBBF0000FBBF0000;
defparam \cp_ready~2 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~3 (
	.dataa(!mem_used_1),
	.datab(!WideOr0),
	.datac(!waitrequest_reset_override),
	.datad(!wait_latency_counter_1),
	.datae(!wait_latency_counter_0),
	.dataf(!\local_write~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready2),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~3 .extended_lut = "off";
defparam \cp_ready~3 .lut_mask = 64'h00000F0002000D00;
defparam \cp_ready~3 .shared_arith = "off";

cyclonev_lcell_comb \rf_source_valid~0 (
	.dataa(!in_data_reg_68),
	.datab(!out_valid_reg),
	.datac(!nxt_out_eop),
	.datad(!in_data_reg_69),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rf_source_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_source_valid~0 .extended_lut = "off";
defparam \rf_source_valid~0 .lut_mask = 64'h0133013301330133;
defparam \rf_source_valid~0 .shared_arith = "off";

cyclonev_lcell_comb local_write(
	.dataa(!in_data_reg_68),
	.datab(!out_valid_reg),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\local_write~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam local_write.extended_lut = "off";
defparam local_write.lut_mask = 64'h1111111111111111;
defparam local_write.shared_arith = "off";

cyclonev_lcell_comb \cp_ready~1 (
	.dataa(!in_narrow_reg),
	.datab(!in_byteen_reg_3),
	.datac(!in_byteen_reg_2),
	.datad(!in_byteen_reg_1),
	.datae(!in_byteen_reg_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cp_ready~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~1 .extended_lut = "off";
defparam \cp_ready~1 .lut_mask = 64'h8000000080000000;
defparam \cp_ready~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_burst_uncompressor_6 (
	mem_66_0,
	comb,
	last_packet_beat,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	last_packet_beat1,
	reset,
	last_packet_beat2,
	WideOr0,
	read,
	sink_ready,
	clk)/* synthesis synthesis_greybox=0 */;
input 	mem_66_0;
input 	comb;
output 	last_packet_beat;
input 	mem_78_0;
input 	mem_77_0;
input 	mem_76_0;
input 	mem_75_0;
input 	mem_74_0;
output 	last_packet_beat1;
input 	reset;
output 	last_packet_beat2;
input 	WideOr0;
input 	read;
output 	sink_ready;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \burst_uncompress_busy~q ;
wire \burst_uncompress_byte_counter~5_combout ;
wire \burst_uncompress_byte_counter[2]~q ;
wire \burst_uncompress_byte_counter~4_combout ;
wire \burst_uncompress_byte_counter[3]~q ;
wire \Add0~2_combout ;
wire \burst_uncompress_byte_counter~3_combout ;
wire \burst_uncompress_byte_counter[4]~q ;
wire \last_packet_beat~3_combout ;
wire \Add1~0_combout ;
wire \burst_uncompress_byte_counter~6_combout ;
wire \burst_uncompress_byte_counter[7]~q ;
wire \burst_uncompress_byte_counter~0_combout ;
wire \Add0~1_combout ;
wire \Add1~1_combout ;
wire \burst_uncompress_byte_counter~2_combout ;
wire \burst_uncompress_byte_counter[5]~q ;
wire \Add0~0_combout ;
wire \burst_uncompress_byte_counter~1_combout ;
wire \burst_uncompress_byte_counter[6]~q ;


cyclonev_lcell_comb \last_packet_beat~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!\burst_uncompress_byte_counter[5]~q ),
	.datad(!\burst_uncompress_byte_counter[4]~q ),
	.datae(!\burst_uncompress_byte_counter[3]~q ),
	.dataf(!\burst_uncompress_byte_counter[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~0 .extended_lut = "off";
defparam \last_packet_beat~0 .lut_mask = 64'h0000000040000000;
defparam \last_packet_beat~0 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~1 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_78_0),
	.datac(!mem_77_0),
	.datad(!mem_76_0),
	.datae(!mem_75_0),
	.dataf(!mem_74_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat1),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~1 .extended_lut = "off";
defparam \last_packet_beat~1 .lut_mask = 64'h0000000080000000;
defparam \last_packet_beat~1 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~2 (
	.dataa(!comb),
	.datab(!mem_66_0),
	.datac(!last_packet_beat),
	.datad(!last_packet_beat1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat2),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~2 .extended_lut = "off";
defparam \last_packet_beat~2 .lut_mask = 64'h3222322232223222;
defparam \last_packet_beat~2 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!comb),
	.datad(!last_packet_beat2),
	.datae(!WideOr0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~0 .extended_lut = "off";
defparam \sink_ready~0 .lut_mask = 64'h00000F0000000F00;
defparam \sink_ready~0 .shared_arith = "off";

dffeas burst_uncompress_busy(
	.clk(clk),
	.d(last_packet_beat2),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_busy~q ),
	.prn(vcc));
defparam burst_uncompress_busy.is_wysiwyg = "true";
defparam burst_uncompress_busy.power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~5 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_74_0),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(!last_packet_beat2),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~5 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~5 .lut_mask = 64'h00C800FA00C800FA;
defparam \burst_uncompress_byte_counter~5 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[2] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[2]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[2] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[2] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~4 (
	.dataa(!mem_75_0),
	.datab(!mem_74_0),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(!last_packet_beat2),
	.dataf(!\burst_uncompress_byte_counter~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~4 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~4 .lut_mask = 64'h000099990000F00F;
defparam \burst_uncompress_byte_counter~4 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[3] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[3]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[3] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[3] .power_up = "low";

cyclonev_lcell_comb \Add0~2 (
	.dataa(!\burst_uncompress_byte_counter[4]~q ),
	.datab(!\burst_uncompress_byte_counter[3]~q ),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~2 .extended_lut = "off";
defparam \Add0~2 .lut_mask = 64'h6A6A6A6A6A6A6A6A;
defparam \Add0~2 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~3 (
	.dataa(!mem_76_0),
	.datab(!mem_75_0),
	.datac(!mem_74_0),
	.datad(!last_packet_beat2),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add0~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~3 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~3 .lut_mask = 64'h009500FF00950000;
defparam \burst_uncompress_byte_counter~3 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[4] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[4]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[4] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[4] .power_up = "low";

cyclonev_lcell_comb \last_packet_beat~3 (
	.dataa(!\burst_uncompress_byte_counter[6]~q ),
	.datab(!\burst_uncompress_byte_counter[5]~q ),
	.datac(!\burst_uncompress_byte_counter[4]~q ),
	.datad(!\burst_uncompress_byte_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_packet_beat~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~3 .extended_lut = "off";
defparam \last_packet_beat~3 .lut_mask = 64'h8000800080008000;
defparam \last_packet_beat~3 .shared_arith = "off";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!mem_77_0),
	.datab(!mem_76_0),
	.datac(!mem_75_0),
	.datad(!mem_74_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h8000800080008000;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~6 (
	.dataa(!mem_78_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat2),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~6 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~6 .lut_mask = 64'h0000000C0A0A000C;
defparam \burst_uncompress_byte_counter~6 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[7] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[7]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[7] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[7] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[2]~q ),
	.datac(!\last_packet_beat~3_combout ),
	.datad(!\burst_uncompress_byte_counter[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~0 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~0 .lut_mask = 64'h5155515551555155;
defparam \burst_uncompress_byte_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!mem_77_0),
	.datab(!mem_76_0),
	.datac(!mem_75_0),
	.datad(!mem_74_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~2 (
	.dataa(!last_packet_beat2),
	.datab(!\burst_uncompress_byte_counter~0_combout ),
	.datac(!\Add0~1_combout ),
	.datad(!\Add1~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~2 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~2 .lut_mask = 64'h5410541054105410;
defparam \burst_uncompress_byte_counter~2 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[5] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[5]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[5] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[5] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h8000800080008000;
defparam \Add0~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~1 (
	.dataa(!mem_78_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat2),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~1 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~1 .lut_mask = 64'h0505030C0A0A030C;
defparam \burst_uncompress_byte_counter~1 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[6] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[6]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[6] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[6] .power_up = "low";

endmodule

module spw_babasu_altera_merlin_slave_agent_7 (
	waitrequest_reset_override,
	stateST_COMP_TRANS,
	out_valid_reg,
	mem_used_1,
	in_narrow_reg,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	WideOr0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	in_data_reg_68,
	cp_ready,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_129_0,
	mem_used_01,
	mem_66_0,
	comb,
	last_packet_beat,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	last_packet_beat1,
	altera_reset_synchronizer_int_chain_out,
	m0_write1,
	nxt_out_eop,
	cp_ready1,
	last_packet_beat2,
	WideOr01,
	read,
	cp_ready2,
	in_data_reg_69,
	rf_source_valid,
	rf_sink_ready,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	waitrequest_reset_override;
input 	stateST_COMP_TRANS;
input 	out_valid_reg;
input 	mem_used_1;
input 	in_narrow_reg;
input 	in_byteen_reg_3;
input 	in_byteen_reg_2;
input 	in_byteen_reg_1;
input 	in_byteen_reg_0;
output 	WideOr0;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	in_data_reg_68;
output 	cp_ready;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	mem_129_0;
input 	mem_used_01;
input 	mem_66_0;
output 	comb;
output 	last_packet_beat;
input 	mem_78_0;
input 	mem_77_0;
input 	mem_76_0;
input 	mem_75_0;
input 	mem_74_0;
output 	last_packet_beat1;
input 	altera_reset_synchronizer_int_chain_out;
output 	m0_write1;
input 	nxt_out_eop;
output 	cp_ready1;
output 	last_packet_beat2;
input 	WideOr01;
input 	read;
output 	cp_ready2;
input 	in_data_reg_69;
output 	rf_source_valid;
output 	rf_sink_ready;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \local_write~combout ;
wire \cp_ready~1_combout ;
wire \cp_ready~2_combout ;


spw_babasu_altera_merlin_burst_uncompressor_7 uncompressor(
	.mem_66_0(mem_66_0),
	.comb(comb),
	.last_packet_beat(last_packet_beat),
	.mem_78_0(mem_78_0),
	.mem_77_0(mem_77_0),
	.mem_76_0(mem_76_0),
	.mem_75_0(mem_75_0),
	.mem_74_0(mem_74_0),
	.last_packet_beat1(last_packet_beat1),
	.reset(altera_reset_synchronizer_int_chain_out),
	.last_packet_beat2(last_packet_beat2),
	.WideOr0(WideOr01),
	.read(read),
	.sink_ready(rf_sink_ready),
	.clk(clk_clk));

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!in_narrow_reg),
	.datac(!in_byteen_reg_3),
	.datad(!in_byteen_reg_2),
	.datae(!in_byteen_reg_1),
	.dataf(!in_byteen_reg_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h1FFFFFFFFFFFFFFF;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~0 (
	.dataa(!waitrequest_reset_override),
	.datab(!mem_used_1),
	.datac(!WideOr0),
	.datad(!wait_latency_counter_1),
	.datae(!wait_latency_counter_0),
	.dataf(!\local_write~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~0 .extended_lut = "off";
defparam \cp_ready~0 .lut_mask = 64'hC0C0C4C0C4C0C0C0;
defparam \cp_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \comb~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_129_0),
	.datad(!mem_used_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(comb),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~0 .extended_lut = "off";
defparam \comb~0 .lut_mask = 64'h007F007F007F007F;
defparam \comb~0 .shared_arith = "off";

cyclonev_lcell_comb m0_write(
	.dataa(!mem_used_1),
	.datab(!WideOr0),
	.datac(!\local_write~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write1),
	.sumout(),
	.cout(),
	.shareout());
defparam m0_write.extended_lut = "off";
defparam m0_write.lut_mask = 64'h0202020202020202;
defparam m0_write.shared_arith = "off";

cyclonev_lcell_comb \cp_ready~3 (
	.dataa(!mem_used_1),
	.datab(!in_narrow_reg),
	.datac(!\cp_ready~1_combout ),
	.datad(!\cp_ready~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~3 .extended_lut = "off";
defparam \cp_ready~3 .lut_mask = 64'h08AA08AA08AA08AA;
defparam \cp_ready~3 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~4 (
	.dataa(!waitrequest_reset_override),
	.datab(!mem_used_1),
	.datac(!WideOr0),
	.datad(!wait_latency_counter_1),
	.datae(!wait_latency_counter_0),
	.dataf(!\local_write~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready2),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~4 .extended_lut = "off";
defparam \cp_ready~4 .lut_mask = 64'h0000550004005100;
defparam \cp_ready~4 .shared_arith = "off";

cyclonev_lcell_comb \rf_source_valid~0 (
	.dataa(!in_data_reg_68),
	.datab(!out_valid_reg),
	.datac(!nxt_out_eop),
	.datad(!in_data_reg_69),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rf_source_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_source_valid~0 .extended_lut = "off";
defparam \rf_source_valid~0 .lut_mask = 64'h0133013301330133;
defparam \rf_source_valid~0 .shared_arith = "off";

cyclonev_lcell_comb local_write(
	.dataa(!in_data_reg_68),
	.datab(!out_valid_reg),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\local_write~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam local_write.extended_lut = "off";
defparam local_write.lut_mask = 64'h1111111111111111;
defparam local_write.shared_arith = "off";

cyclonev_lcell_comb \cp_ready~1 (
	.dataa(!in_byteen_reg_3),
	.datab(!in_byteen_reg_2),
	.datac(!in_byteen_reg_1),
	.datad(!in_byteen_reg_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cp_ready~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~1 .extended_lut = "off";
defparam \cp_ready~1 .lut_mask = 64'h8000800080008000;
defparam \cp_ready~1 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~2 (
	.dataa(!waitrequest_reset_override),
	.datab(!wait_latency_counter_1),
	.datac(!wait_latency_counter_0),
	.datad(!\local_write~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cp_ready~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~2 .extended_lut = "off";
defparam \cp_ready~2 .lut_mask = 64'h0440044004400440;
defparam \cp_ready~2 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_burst_uncompressor_7 (
	mem_66_0,
	comb,
	last_packet_beat,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	last_packet_beat1,
	reset,
	last_packet_beat2,
	WideOr0,
	read,
	sink_ready,
	clk)/* synthesis synthesis_greybox=0 */;
input 	mem_66_0;
input 	comb;
output 	last_packet_beat;
input 	mem_78_0;
input 	mem_77_0;
input 	mem_76_0;
input 	mem_75_0;
input 	mem_74_0;
output 	last_packet_beat1;
input 	reset;
output 	last_packet_beat2;
input 	WideOr0;
input 	read;
output 	sink_ready;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \burst_uncompress_busy~q ;
wire \burst_uncompress_byte_counter~5_combout ;
wire \burst_uncompress_byte_counter[2]~q ;
wire \burst_uncompress_byte_counter~4_combout ;
wire \burst_uncompress_byte_counter[3]~q ;
wire \Add0~2_combout ;
wire \burst_uncompress_byte_counter~3_combout ;
wire \burst_uncompress_byte_counter[4]~q ;
wire \last_packet_beat~3_combout ;
wire \Add1~0_combout ;
wire \burst_uncompress_byte_counter~6_combout ;
wire \burst_uncompress_byte_counter[7]~q ;
wire \burst_uncompress_byte_counter~0_combout ;
wire \Add0~1_combout ;
wire \Add1~1_combout ;
wire \burst_uncompress_byte_counter~2_combout ;
wire \burst_uncompress_byte_counter[5]~q ;
wire \Add0~0_combout ;
wire \burst_uncompress_byte_counter~1_combout ;
wire \burst_uncompress_byte_counter[6]~q ;


cyclonev_lcell_comb \last_packet_beat~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!\burst_uncompress_byte_counter[5]~q ),
	.datad(!\burst_uncompress_byte_counter[4]~q ),
	.datae(!\burst_uncompress_byte_counter[3]~q ),
	.dataf(!\burst_uncompress_byte_counter[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~0 .extended_lut = "off";
defparam \last_packet_beat~0 .lut_mask = 64'h0000000040000000;
defparam \last_packet_beat~0 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~1 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_78_0),
	.datac(!mem_77_0),
	.datad(!mem_76_0),
	.datae(!mem_75_0),
	.dataf(!mem_74_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat1),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~1 .extended_lut = "off";
defparam \last_packet_beat~1 .lut_mask = 64'h0000000080000000;
defparam \last_packet_beat~1 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~2 (
	.dataa(!comb),
	.datab(!mem_66_0),
	.datac(!last_packet_beat),
	.datad(!last_packet_beat1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat2),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~2 .extended_lut = "off";
defparam \last_packet_beat~2 .lut_mask = 64'h3222322232223222;
defparam \last_packet_beat~2 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!comb),
	.datad(!last_packet_beat2),
	.datae(!WideOr0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~0 .extended_lut = "off";
defparam \sink_ready~0 .lut_mask = 64'h00000F0000000F00;
defparam \sink_ready~0 .shared_arith = "off";

dffeas burst_uncompress_busy(
	.clk(clk),
	.d(last_packet_beat2),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_busy~q ),
	.prn(vcc));
defparam burst_uncompress_busy.is_wysiwyg = "true";
defparam burst_uncompress_busy.power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~5 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_74_0),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(!last_packet_beat2),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~5 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~5 .lut_mask = 64'h00C800FA00C800FA;
defparam \burst_uncompress_byte_counter~5 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[2] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[2]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[2] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[2] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~4 (
	.dataa(!mem_75_0),
	.datab(!mem_74_0),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(!last_packet_beat2),
	.dataf(!\burst_uncompress_byte_counter~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~4 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~4 .lut_mask = 64'h000099990000F00F;
defparam \burst_uncompress_byte_counter~4 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[3] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[3]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[3] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[3] .power_up = "low";

cyclonev_lcell_comb \Add0~2 (
	.dataa(!\burst_uncompress_byte_counter[4]~q ),
	.datab(!\burst_uncompress_byte_counter[3]~q ),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~2 .extended_lut = "off";
defparam \Add0~2 .lut_mask = 64'h6A6A6A6A6A6A6A6A;
defparam \Add0~2 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~3 (
	.dataa(!mem_76_0),
	.datab(!mem_75_0),
	.datac(!mem_74_0),
	.datad(!last_packet_beat2),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add0~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~3 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~3 .lut_mask = 64'h009500FF00950000;
defparam \burst_uncompress_byte_counter~3 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[4] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[4]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[4] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[4] .power_up = "low";

cyclonev_lcell_comb \last_packet_beat~3 (
	.dataa(!\burst_uncompress_byte_counter[6]~q ),
	.datab(!\burst_uncompress_byte_counter[5]~q ),
	.datac(!\burst_uncompress_byte_counter[4]~q ),
	.datad(!\burst_uncompress_byte_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_packet_beat~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~3 .extended_lut = "off";
defparam \last_packet_beat~3 .lut_mask = 64'h8000800080008000;
defparam \last_packet_beat~3 .shared_arith = "off";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!mem_77_0),
	.datab(!mem_76_0),
	.datac(!mem_75_0),
	.datad(!mem_74_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h8000800080008000;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~6 (
	.dataa(!mem_78_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat2),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~6 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~6 .lut_mask = 64'h0000000C0A0A000C;
defparam \burst_uncompress_byte_counter~6 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[7] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[7]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[7] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[7] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[2]~q ),
	.datac(!\last_packet_beat~3_combout ),
	.datad(!\burst_uncompress_byte_counter[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~0 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~0 .lut_mask = 64'h5155515551555155;
defparam \burst_uncompress_byte_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!mem_77_0),
	.datab(!mem_76_0),
	.datac(!mem_75_0),
	.datad(!mem_74_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~2 (
	.dataa(!last_packet_beat2),
	.datab(!\burst_uncompress_byte_counter~0_combout ),
	.datac(!\Add0~1_combout ),
	.datad(!\Add1~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~2 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~2 .lut_mask = 64'h5410541054105410;
defparam \burst_uncompress_byte_counter~2 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[5] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[5]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[5] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[5] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h8000800080008000;
defparam \Add0~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~1 (
	.dataa(!mem_78_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat2),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~1 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~1 .lut_mask = 64'h0505030C0A0A030C;
defparam \burst_uncompress_byte_counter~1 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[6] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[6]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[6] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[6] .power_up = "low";

endmodule

module spw_babasu_altera_merlin_slave_agent_8 (
	h2f_RREADY_0,
	waitrequest_reset_override,
	stateST_COMP_TRANS,
	mem_used_1,
	in_data_reg_69,
	in_narrow_reg,
	wait_latency_counter_1,
	wait_latency_counter_0,
	cp_ready,
	cp_ready1,
	empty,
	mem_66_0,
	mem_used_0,
	last_packet_beat,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	last_packet_beat1,
	altera_reset_synchronizer_int_chain_out,
	last_packet_beat2,
	cp_ready2,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_RREADY_0;
input 	waitrequest_reset_override;
input 	stateST_COMP_TRANS;
input 	mem_used_1;
input 	in_data_reg_69;
input 	in_narrow_reg;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
output 	cp_ready;
output 	cp_ready1;
input 	empty;
input 	mem_66_0;
input 	mem_used_0;
output 	last_packet_beat;
input 	mem_78_0;
input 	mem_77_0;
input 	mem_76_0;
input 	mem_75_0;
input 	mem_74_0;
output 	last_packet_beat1;
input 	altera_reset_synchronizer_int_chain_out;
output 	last_packet_beat2;
output 	cp_ready2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



spw_babasu_altera_merlin_burst_uncompressor_8 uncompressor(
	.h2f_RREADY_0(h2f_RREADY_0),
	.empty(empty),
	.mem_66_0(mem_66_0),
	.mem_used_0(mem_used_0),
	.last_packet_beat(last_packet_beat),
	.mem_78_0(mem_78_0),
	.mem_77_0(mem_77_0),
	.mem_76_0(mem_76_0),
	.mem_75_0(mem_75_0),
	.mem_74_0(mem_74_0),
	.last_packet_beat1(last_packet_beat1),
	.reset(altera_reset_synchronizer_int_chain_out),
	.last_packet_beat2(last_packet_beat2),
	.clk(clk_clk));

cyclonev_lcell_comb \cp_ready~0 (
	.dataa(!waitrequest_reset_override),
	.datab(!in_data_reg_69),
	.datac(!stateST_COMP_TRANS),
	.datad(!in_narrow_reg),
	.datae(!wait_latency_counter_1),
	.dataf(!wait_latency_counter_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~0 .extended_lut = "off";
defparam \cp_ready~0 .lut_mask = 64'hCCC0CCC0DDD5CCC0;
defparam \cp_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~1 (
	.dataa(!mem_used_1),
	.datab(!cp_ready),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~1 .extended_lut = "off";
defparam \cp_ready~1 .lut_mask = 64'h2222222222222222;
defparam \cp_ready~1 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~2 (
	.dataa(!waitrequest_reset_override),
	.datab(!in_data_reg_69),
	.datac(!in_narrow_reg),
	.datad(!wait_latency_counter_1),
	.datae(!wait_latency_counter_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready2),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~2 .extended_lut = "off";
defparam \cp_ready~2 .lut_mask = 64'hC0C0D5C0C0C0D5C0;
defparam \cp_ready~2 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_burst_uncompressor_8 (
	h2f_RREADY_0,
	empty,
	mem_66_0,
	mem_used_0,
	last_packet_beat,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	last_packet_beat1,
	reset,
	last_packet_beat2,
	clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_RREADY_0;
input 	empty;
input 	mem_66_0;
input 	mem_used_0;
output 	last_packet_beat;
input 	mem_78_0;
input 	mem_77_0;
input 	mem_76_0;
input 	mem_75_0;
input 	mem_74_0;
output 	last_packet_beat1;
input 	reset;
output 	last_packet_beat2;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always0~0_combout ;
wire \burst_uncompress_busy~q ;
wire \burst_uncompress_byte_counter~5_combout ;
wire \burst_uncompress_byte_counter[2]~q ;
wire \burst_uncompress_byte_counter~4_combout ;
wire \burst_uncompress_byte_counter[3]~q ;
wire \Add0~2_combout ;
wire \burst_uncompress_byte_counter~3_combout ;
wire \burst_uncompress_byte_counter[4]~q ;
wire \last_packet_beat~3_combout ;
wire \Add1~0_combout ;
wire \burst_uncompress_byte_counter~6_combout ;
wire \burst_uncompress_byte_counter[7]~q ;
wire \burst_uncompress_byte_counter~0_combout ;
wire \Add0~1_combout ;
wire \Add1~1_combout ;
wire \burst_uncompress_byte_counter~2_combout ;
wire \burst_uncompress_byte_counter[5]~q ;
wire \Add0~0_combout ;
wire \burst_uncompress_byte_counter~1_combout ;
wire \burst_uncompress_byte_counter[6]~q ;


cyclonev_lcell_comb \last_packet_beat~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!\burst_uncompress_byte_counter[5]~q ),
	.datad(!\burst_uncompress_byte_counter[4]~q ),
	.datae(!\burst_uncompress_byte_counter[3]~q ),
	.dataf(!\burst_uncompress_byte_counter[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~0 .extended_lut = "off";
defparam \last_packet_beat~0 .lut_mask = 64'h0000000040000000;
defparam \last_packet_beat~0 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~1 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_78_0),
	.datac(!mem_77_0),
	.datad(!mem_76_0),
	.datae(!mem_75_0),
	.dataf(!mem_74_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat1),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~1 .extended_lut = "off";
defparam \last_packet_beat~1 .lut_mask = 64'h0000000080000000;
defparam \last_packet_beat~1 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~2 (
	.dataa(!empty),
	.datab(!mem_66_0),
	.datac(!mem_used_0),
	.datad(!last_packet_beat),
	.datae(!last_packet_beat1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat2),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~2 .extended_lut = "off";
defparam \last_packet_beat~2 .lut_mask = 64'h3331313133313131;
defparam \last_packet_beat~2 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!h2f_RREADY_0),
	.datab(!empty),
	.datac(!mem_used_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'h0404040404040404;
defparam \always0~0 .shared_arith = "off";

dffeas burst_uncompress_busy(
	.clk(clk),
	.d(last_packet_beat2),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_busy~q ),
	.prn(vcc));
defparam burst_uncompress_busy.is_wysiwyg = "true";
defparam burst_uncompress_busy.power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~5 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_74_0),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(!last_packet_beat2),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~5 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~5 .lut_mask = 64'h00C800FA00C800FA;
defparam \burst_uncompress_byte_counter~5 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[2] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[2]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[2] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[2] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~4 (
	.dataa(!mem_75_0),
	.datab(!mem_74_0),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(!last_packet_beat2),
	.dataf(!\burst_uncompress_byte_counter~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~4 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~4 .lut_mask = 64'h000099990000F00F;
defparam \burst_uncompress_byte_counter~4 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[3] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[3]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[3] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[3] .power_up = "low";

cyclonev_lcell_comb \Add0~2 (
	.dataa(!\burst_uncompress_byte_counter[4]~q ),
	.datab(!\burst_uncompress_byte_counter[3]~q ),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~2 .extended_lut = "off";
defparam \Add0~2 .lut_mask = 64'h6A6A6A6A6A6A6A6A;
defparam \Add0~2 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~3 (
	.dataa(!mem_76_0),
	.datab(!mem_75_0),
	.datac(!mem_74_0),
	.datad(!last_packet_beat2),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add0~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~3 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~3 .lut_mask = 64'h009500FF00950000;
defparam \burst_uncompress_byte_counter~3 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[4] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[4]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[4] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[4] .power_up = "low";

cyclonev_lcell_comb \last_packet_beat~3 (
	.dataa(!\burst_uncompress_byte_counter[6]~q ),
	.datab(!\burst_uncompress_byte_counter[5]~q ),
	.datac(!\burst_uncompress_byte_counter[4]~q ),
	.datad(!\burst_uncompress_byte_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_packet_beat~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~3 .extended_lut = "off";
defparam \last_packet_beat~3 .lut_mask = 64'h8000800080008000;
defparam \last_packet_beat~3 .shared_arith = "off";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!mem_77_0),
	.datab(!mem_76_0),
	.datac(!mem_75_0),
	.datad(!mem_74_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h8000800080008000;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~6 (
	.dataa(!mem_78_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat2),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~6 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~6 .lut_mask = 64'h0000000C0A0A000C;
defparam \burst_uncompress_byte_counter~6 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[7] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[7]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[7] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[7] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[2]~q ),
	.datac(!\last_packet_beat~3_combout ),
	.datad(!\burst_uncompress_byte_counter[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~0 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~0 .lut_mask = 64'h5155515551555155;
defparam \burst_uncompress_byte_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!mem_77_0),
	.datab(!mem_76_0),
	.datac(!mem_75_0),
	.datad(!mem_74_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~2 (
	.dataa(!last_packet_beat2),
	.datab(!\burst_uncompress_byte_counter~0_combout ),
	.datac(!\Add0~1_combout ),
	.datad(!\Add1~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~2 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~2 .lut_mask = 64'h5410541054105410;
defparam \burst_uncompress_byte_counter~2 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[5] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[5]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[5] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[5] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h8000800080008000;
defparam \Add0~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~1 (
	.dataa(!mem_78_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat2),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~1 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~1 .lut_mask = 64'h0505030C0A0A030C;
defparam \burst_uncompress_byte_counter~1 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[6] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[6]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[6] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[6] .power_up = "low";

endmodule

module spw_babasu_altera_merlin_slave_agent_9 (
	waitrequest_reset_override,
	stateST_COMP_TRANS,
	out_valid_reg,
	mem_used_1,
	in_narrow_reg,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	WideOr0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	in_data_reg_68,
	cp_ready,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_129_0,
	mem_used_01,
	mem_66_0,
	comb,
	last_packet_beat,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	last_packet_beat1,
	altera_reset_synchronizer_int_chain_out,
	m0_write1,
	nxt_out_eop,
	cp_ready1,
	cp_ready2,
	last_packet_beat2,
	WideOr01,
	read,
	cp_ready3,
	in_data_reg_69,
	rf_source_valid,
	rf_sink_ready,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	waitrequest_reset_override;
input 	stateST_COMP_TRANS;
input 	out_valid_reg;
input 	mem_used_1;
input 	in_narrow_reg;
input 	in_byteen_reg_3;
input 	in_byteen_reg_2;
input 	in_byteen_reg_1;
input 	in_byteen_reg_0;
output 	WideOr0;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	in_data_reg_68;
output 	cp_ready;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	mem_129_0;
input 	mem_used_01;
input 	mem_66_0;
output 	comb;
output 	last_packet_beat;
input 	mem_78_0;
input 	mem_77_0;
input 	mem_76_0;
input 	mem_75_0;
input 	mem_74_0;
output 	last_packet_beat1;
input 	altera_reset_synchronizer_int_chain_out;
output 	m0_write1;
input 	nxt_out_eop;
output 	cp_ready1;
output 	cp_ready2;
output 	last_packet_beat2;
input 	WideOr01;
input 	read;
output 	cp_ready3;
input 	in_data_reg_69;
output 	rf_source_valid;
output 	rf_sink_ready;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \local_write~combout ;


spw_babasu_altera_merlin_burst_uncompressor_9 uncompressor(
	.mem_66_0(mem_66_0),
	.comb(comb),
	.last_packet_beat(last_packet_beat),
	.mem_78_0(mem_78_0),
	.mem_77_0(mem_77_0),
	.mem_76_0(mem_76_0),
	.mem_75_0(mem_75_0),
	.mem_74_0(mem_74_0),
	.last_packet_beat1(last_packet_beat1),
	.reset(altera_reset_synchronizer_int_chain_out),
	.last_packet_beat2(last_packet_beat2),
	.WideOr0(WideOr01),
	.read(read),
	.sink_ready(rf_sink_ready),
	.clk(clk_clk));

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!in_narrow_reg),
	.datac(!in_byteen_reg_3),
	.datad(!in_byteen_reg_2),
	.datae(!in_byteen_reg_1),
	.dataf(!in_byteen_reg_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h1FFFFFFFFFFFFFFF;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~0 (
	.dataa(!waitrequest_reset_override),
	.datab(!mem_used_1),
	.datac(!WideOr0),
	.datad(!wait_latency_counter_1),
	.datae(!wait_latency_counter_0),
	.dataf(!\local_write~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~0 .extended_lut = "off";
defparam \cp_ready~0 .lut_mask = 64'hC0C0C4C0C4C0C0C0;
defparam \cp_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \comb~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_129_0),
	.datad(!mem_used_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(comb),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~0 .extended_lut = "off";
defparam \comb~0 .lut_mask = 64'h007F007F007F007F;
defparam \comb~0 .shared_arith = "off";

cyclonev_lcell_comb m0_write(
	.dataa(!mem_used_1),
	.datab(!WideOr0),
	.datac(!\local_write~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write1),
	.sumout(),
	.cout(),
	.shareout());
defparam m0_write.extended_lut = "off";
defparam m0_write.lut_mask = 64'h0202020202020202;
defparam m0_write.shared_arith = "off";

cyclonev_lcell_comb \cp_ready~1 (
	.dataa(!in_narrow_reg),
	.datab(!in_byteen_reg_3),
	.datac(!in_byteen_reg_2),
	.datad(!in_byteen_reg_1),
	.datae(!in_byteen_reg_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~1 .extended_lut = "off";
defparam \cp_ready~1 .lut_mask = 64'h8000000080000000;
defparam \cp_ready~1 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~2 (
	.dataa(!waitrequest_reset_override),
	.datab(!wait_latency_counter_1),
	.datac(!wait_latency_counter_0),
	.datad(!\local_write~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready2),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~2 .extended_lut = "off";
defparam \cp_ready~2 .lut_mask = 64'h0440044004400440;
defparam \cp_ready~2 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~3 (
	.dataa(!waitrequest_reset_override),
	.datab(!mem_used_1),
	.datac(!WideOr0),
	.datad(!wait_latency_counter_1),
	.datae(!wait_latency_counter_0),
	.dataf(!\local_write~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready3),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~3 .extended_lut = "off";
defparam \cp_ready~3 .lut_mask = 64'h0000550004005100;
defparam \cp_ready~3 .shared_arith = "off";

cyclonev_lcell_comb \rf_source_valid~0 (
	.dataa(!in_data_reg_68),
	.datab(!out_valid_reg),
	.datac(!nxt_out_eop),
	.datad(!in_data_reg_69),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rf_source_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_source_valid~0 .extended_lut = "off";
defparam \rf_source_valid~0 .lut_mask = 64'h0133013301330133;
defparam \rf_source_valid~0 .shared_arith = "off";

cyclonev_lcell_comb local_write(
	.dataa(!in_data_reg_68),
	.datab(!out_valid_reg),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\local_write~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam local_write.extended_lut = "off";
defparam local_write.lut_mask = 64'h1111111111111111;
defparam local_write.shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_burst_uncompressor_9 (
	mem_66_0,
	comb,
	last_packet_beat,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	last_packet_beat1,
	reset,
	last_packet_beat2,
	WideOr0,
	read,
	sink_ready,
	clk)/* synthesis synthesis_greybox=0 */;
input 	mem_66_0;
input 	comb;
output 	last_packet_beat;
input 	mem_78_0;
input 	mem_77_0;
input 	mem_76_0;
input 	mem_75_0;
input 	mem_74_0;
output 	last_packet_beat1;
input 	reset;
output 	last_packet_beat2;
input 	WideOr0;
input 	read;
output 	sink_ready;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \burst_uncompress_busy~q ;
wire \burst_uncompress_byte_counter~5_combout ;
wire \burst_uncompress_byte_counter[2]~q ;
wire \burst_uncompress_byte_counter~4_combout ;
wire \burst_uncompress_byte_counter[3]~q ;
wire \Add0~2_combout ;
wire \burst_uncompress_byte_counter~3_combout ;
wire \burst_uncompress_byte_counter[4]~q ;
wire \last_packet_beat~3_combout ;
wire \Add1~0_combout ;
wire \burst_uncompress_byte_counter~6_combout ;
wire \burst_uncompress_byte_counter[7]~q ;
wire \burst_uncompress_byte_counter~0_combout ;
wire \Add0~1_combout ;
wire \Add1~1_combout ;
wire \burst_uncompress_byte_counter~2_combout ;
wire \burst_uncompress_byte_counter[5]~q ;
wire \Add0~0_combout ;
wire \burst_uncompress_byte_counter~1_combout ;
wire \burst_uncompress_byte_counter[6]~q ;


cyclonev_lcell_comb \last_packet_beat~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!\burst_uncompress_byte_counter[5]~q ),
	.datad(!\burst_uncompress_byte_counter[4]~q ),
	.datae(!\burst_uncompress_byte_counter[3]~q ),
	.dataf(!\burst_uncompress_byte_counter[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~0 .extended_lut = "off";
defparam \last_packet_beat~0 .lut_mask = 64'h0000000040000000;
defparam \last_packet_beat~0 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~1 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_78_0),
	.datac(!mem_77_0),
	.datad(!mem_76_0),
	.datae(!mem_75_0),
	.dataf(!mem_74_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat1),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~1 .extended_lut = "off";
defparam \last_packet_beat~1 .lut_mask = 64'h0000000080000000;
defparam \last_packet_beat~1 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~2 (
	.dataa(!comb),
	.datab(!mem_66_0),
	.datac(!last_packet_beat),
	.datad(!last_packet_beat1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat2),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~2 .extended_lut = "off";
defparam \last_packet_beat~2 .lut_mask = 64'h3222322232223222;
defparam \last_packet_beat~2 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!comb),
	.datad(!last_packet_beat2),
	.datae(!WideOr0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~0 .extended_lut = "off";
defparam \sink_ready~0 .lut_mask = 64'h00000F0000000F00;
defparam \sink_ready~0 .shared_arith = "off";

dffeas burst_uncompress_busy(
	.clk(clk),
	.d(last_packet_beat2),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_busy~q ),
	.prn(vcc));
defparam burst_uncompress_busy.is_wysiwyg = "true";
defparam burst_uncompress_busy.power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~5 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_74_0),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(!last_packet_beat2),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~5 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~5 .lut_mask = 64'h00C800FA00C800FA;
defparam \burst_uncompress_byte_counter~5 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[2] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[2]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[2] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[2] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~4 (
	.dataa(!mem_75_0),
	.datab(!mem_74_0),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(!last_packet_beat2),
	.dataf(!\burst_uncompress_byte_counter~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~4 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~4 .lut_mask = 64'h000099990000F00F;
defparam \burst_uncompress_byte_counter~4 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[3] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[3]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[3] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[3] .power_up = "low";

cyclonev_lcell_comb \Add0~2 (
	.dataa(!\burst_uncompress_byte_counter[4]~q ),
	.datab(!\burst_uncompress_byte_counter[3]~q ),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~2 .extended_lut = "off";
defparam \Add0~2 .lut_mask = 64'h6A6A6A6A6A6A6A6A;
defparam \Add0~2 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~3 (
	.dataa(!mem_76_0),
	.datab(!mem_75_0),
	.datac(!mem_74_0),
	.datad(!last_packet_beat2),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add0~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~3 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~3 .lut_mask = 64'h009500FF00950000;
defparam \burst_uncompress_byte_counter~3 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[4] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[4]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[4] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[4] .power_up = "low";

cyclonev_lcell_comb \last_packet_beat~3 (
	.dataa(!\burst_uncompress_byte_counter[6]~q ),
	.datab(!\burst_uncompress_byte_counter[5]~q ),
	.datac(!\burst_uncompress_byte_counter[4]~q ),
	.datad(!\burst_uncompress_byte_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_packet_beat~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~3 .extended_lut = "off";
defparam \last_packet_beat~3 .lut_mask = 64'h8000800080008000;
defparam \last_packet_beat~3 .shared_arith = "off";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!mem_77_0),
	.datab(!mem_76_0),
	.datac(!mem_75_0),
	.datad(!mem_74_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h8000800080008000;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~6 (
	.dataa(!mem_78_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat2),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~6 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~6 .lut_mask = 64'h0000000C0A0A000C;
defparam \burst_uncompress_byte_counter~6 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[7] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[7]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[7] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[7] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[2]~q ),
	.datac(!\last_packet_beat~3_combout ),
	.datad(!\burst_uncompress_byte_counter[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~0 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~0 .lut_mask = 64'h5155515551555155;
defparam \burst_uncompress_byte_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!mem_77_0),
	.datab(!mem_76_0),
	.datac(!mem_75_0),
	.datad(!mem_74_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~2 (
	.dataa(!last_packet_beat2),
	.datab(!\burst_uncompress_byte_counter~0_combout ),
	.datac(!\Add0~1_combout ),
	.datad(!\Add1~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~2 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~2 .lut_mask = 64'h5410541054105410;
defparam \burst_uncompress_byte_counter~2 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[5] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[5]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[5] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[5] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h8000800080008000;
defparam \Add0~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~1 (
	.dataa(!mem_78_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat2),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~1 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~1 .lut_mask = 64'h0505030C0A0A030C;
defparam \burst_uncompress_byte_counter~1 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[6] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[6]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[6] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[6] .power_up = "low";

endmodule

module spw_babasu_altera_merlin_slave_agent_10 (
	waitrequest_reset_override,
	stateST_COMP_TRANS,
	out_valid_reg,
	mem_used_1,
	in_narrow_reg,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	WideOr0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	in_data_reg_68,
	cp_ready,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_129_0,
	mem_used_01,
	mem_66_0,
	comb,
	last_packet_beat,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	last_packet_beat1,
	altera_reset_synchronizer_int_chain_out,
	m0_write1,
	nxt_out_eop,
	cp_ready1,
	last_packet_beat2,
	read,
	cp_ready2,
	in_data_reg_69,
	rf_source_valid,
	rp_valid1,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	waitrequest_reset_override;
input 	stateST_COMP_TRANS;
input 	out_valid_reg;
input 	mem_used_1;
input 	in_narrow_reg;
input 	in_byteen_reg_3;
input 	in_byteen_reg_2;
input 	in_byteen_reg_1;
input 	in_byteen_reg_0;
output 	WideOr0;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	in_data_reg_68;
output 	cp_ready;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	mem_129_0;
input 	mem_used_01;
input 	mem_66_0;
output 	comb;
output 	last_packet_beat;
input 	mem_78_0;
input 	mem_77_0;
input 	mem_76_0;
input 	mem_75_0;
input 	mem_74_0;
output 	last_packet_beat1;
input 	altera_reset_synchronizer_int_chain_out;
output 	m0_write1;
input 	nxt_out_eop;
output 	cp_ready1;
output 	last_packet_beat2;
input 	read;
output 	cp_ready2;
input 	in_data_reg_69;
output 	rf_source_valid;
output 	rp_valid1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \local_write~combout ;
wire \cp_ready~1_combout ;
wire \cp_ready~2_combout ;


spw_babasu_altera_merlin_burst_uncompressor_10 uncompressor(
	.mem_66_0(mem_66_0),
	.comb(comb),
	.last_packet_beat(last_packet_beat),
	.mem_78_0(mem_78_0),
	.mem_77_0(mem_77_0),
	.mem_76_0(mem_76_0),
	.mem_75_0(mem_75_0),
	.mem_74_0(mem_74_0),
	.last_packet_beat1(last_packet_beat1),
	.reset(altera_reset_synchronizer_int_chain_out),
	.last_packet_beat2(last_packet_beat2),
	.read(read),
	.clk(clk_clk));

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!in_narrow_reg),
	.datac(!in_byteen_reg_3),
	.datad(!in_byteen_reg_2),
	.datae(!in_byteen_reg_1),
	.dataf(!in_byteen_reg_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h1FFFFFFFFFFFFFFF;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~0 (
	.dataa(!waitrequest_reset_override),
	.datab(!mem_used_1),
	.datac(!WideOr0),
	.datad(!wait_latency_counter_1),
	.datae(!wait_latency_counter_0),
	.dataf(!\local_write~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~0 .extended_lut = "off";
defparam \cp_ready~0 .lut_mask = 64'hC0C0C4C0C4C0C0C0;
defparam \cp_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \comb~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_129_0),
	.datad(!mem_used_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(comb),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~0 .extended_lut = "off";
defparam \comb~0 .lut_mask = 64'h007F007F007F007F;
defparam \comb~0 .shared_arith = "off";

cyclonev_lcell_comb m0_write(
	.dataa(!mem_used_1),
	.datab(!WideOr0),
	.datac(!\local_write~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write1),
	.sumout(),
	.cout(),
	.shareout());
defparam m0_write.extended_lut = "off";
defparam m0_write.lut_mask = 64'h0202020202020202;
defparam m0_write.shared_arith = "off";

cyclonev_lcell_comb \cp_ready~3 (
	.dataa(!mem_used_1),
	.datab(!in_narrow_reg),
	.datac(!\cp_ready~1_combout ),
	.datad(!\cp_ready~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~3 .extended_lut = "off";
defparam \cp_ready~3 .lut_mask = 64'h08AA08AA08AA08AA;
defparam \cp_ready~3 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~4 (
	.dataa(!waitrequest_reset_override),
	.datab(!mem_used_1),
	.datac(!WideOr0),
	.datad(!wait_latency_counter_1),
	.datae(!wait_latency_counter_0),
	.dataf(!\local_write~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready2),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~4 .extended_lut = "off";
defparam \cp_ready~4 .lut_mask = 64'h0000550004005100;
defparam \cp_ready~4 .shared_arith = "off";

cyclonev_lcell_comb \rf_source_valid~0 (
	.dataa(!in_data_reg_68),
	.datab(!out_valid_reg),
	.datac(!nxt_out_eop),
	.datad(!in_data_reg_69),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rf_source_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_source_valid~0 .extended_lut = "off";
defparam \rf_source_valid~0 .lut_mask = 64'h0133013301330133;
defparam \rf_source_valid~0 .shared_arith = "off";

cyclonev_lcell_comb rp_valid(
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_129_0),
	.datad(!mem_used_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rp_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam rp_valid.extended_lut = "off";
defparam rp_valid.lut_mask = 64'h8880888088808880;
defparam rp_valid.shared_arith = "off";

cyclonev_lcell_comb local_write(
	.dataa(!in_data_reg_68),
	.datab(!out_valid_reg),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\local_write~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam local_write.extended_lut = "off";
defparam local_write.lut_mask = 64'h1111111111111111;
defparam local_write.shared_arith = "off";

cyclonev_lcell_comb \cp_ready~1 (
	.dataa(!in_byteen_reg_3),
	.datab(!in_byteen_reg_2),
	.datac(!in_byteen_reg_1),
	.datad(!in_byteen_reg_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cp_ready~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~1 .extended_lut = "off";
defparam \cp_ready~1 .lut_mask = 64'h8000800080008000;
defparam \cp_ready~1 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~2 (
	.dataa(!waitrequest_reset_override),
	.datab(!wait_latency_counter_1),
	.datac(!wait_latency_counter_0),
	.datad(!\local_write~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cp_ready~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~2 .extended_lut = "off";
defparam \cp_ready~2 .lut_mask = 64'h0440044004400440;
defparam \cp_ready~2 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_burst_uncompressor_10 (
	mem_66_0,
	comb,
	last_packet_beat,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	last_packet_beat1,
	reset,
	last_packet_beat2,
	read,
	clk)/* synthesis synthesis_greybox=0 */;
input 	mem_66_0;
input 	comb;
output 	last_packet_beat;
input 	mem_78_0;
input 	mem_77_0;
input 	mem_76_0;
input 	mem_75_0;
input 	mem_74_0;
output 	last_packet_beat1;
input 	reset;
output 	last_packet_beat2;
input 	read;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \burst_uncompress_busy~q ;
wire \burst_uncompress_byte_counter~5_combout ;
wire \burst_uncompress_byte_counter[2]~q ;
wire \burst_uncompress_byte_counter~4_combout ;
wire \burst_uncompress_byte_counter[3]~q ;
wire \Add0~2_combout ;
wire \burst_uncompress_byte_counter~3_combout ;
wire \burst_uncompress_byte_counter[4]~q ;
wire \last_packet_beat~3_combout ;
wire \Add1~0_combout ;
wire \burst_uncompress_byte_counter~6_combout ;
wire \burst_uncompress_byte_counter[7]~q ;
wire \burst_uncompress_byte_counter~0_combout ;
wire \Add0~1_combout ;
wire \Add1~1_combout ;
wire \burst_uncompress_byte_counter~2_combout ;
wire \burst_uncompress_byte_counter[5]~q ;
wire \Add0~0_combout ;
wire \burst_uncompress_byte_counter~1_combout ;
wire \burst_uncompress_byte_counter[6]~q ;


cyclonev_lcell_comb \last_packet_beat~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!\burst_uncompress_byte_counter[5]~q ),
	.datad(!\burst_uncompress_byte_counter[4]~q ),
	.datae(!\burst_uncompress_byte_counter[3]~q ),
	.dataf(!\burst_uncompress_byte_counter[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~0 .extended_lut = "off";
defparam \last_packet_beat~0 .lut_mask = 64'h0000000040000000;
defparam \last_packet_beat~0 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~1 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_78_0),
	.datac(!mem_77_0),
	.datad(!mem_76_0),
	.datae(!mem_75_0),
	.dataf(!mem_74_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat1),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~1 .extended_lut = "off";
defparam \last_packet_beat~1 .lut_mask = 64'h0000000080000000;
defparam \last_packet_beat~1 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~2 (
	.dataa(!comb),
	.datab(!mem_66_0),
	.datac(!last_packet_beat),
	.datad(!last_packet_beat1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat2),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~2 .extended_lut = "off";
defparam \last_packet_beat~2 .lut_mask = 64'h3222322232223222;
defparam \last_packet_beat~2 .shared_arith = "off";

dffeas burst_uncompress_busy(
	.clk(clk),
	.d(last_packet_beat2),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_busy~q ),
	.prn(vcc));
defparam burst_uncompress_busy.is_wysiwyg = "true";
defparam burst_uncompress_busy.power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~5 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_74_0),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(!last_packet_beat2),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~5 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~5 .lut_mask = 64'h00C800FA00C800FA;
defparam \burst_uncompress_byte_counter~5 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[2] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[2]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[2] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[2] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~4 (
	.dataa(!mem_75_0),
	.datab(!mem_74_0),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(!last_packet_beat2),
	.dataf(!\burst_uncompress_byte_counter~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~4 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~4 .lut_mask = 64'h000099990000F00F;
defparam \burst_uncompress_byte_counter~4 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[3] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[3]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[3] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[3] .power_up = "low";

cyclonev_lcell_comb \Add0~2 (
	.dataa(!\burst_uncompress_byte_counter[4]~q ),
	.datab(!\burst_uncompress_byte_counter[3]~q ),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~2 .extended_lut = "off";
defparam \Add0~2 .lut_mask = 64'h6A6A6A6A6A6A6A6A;
defparam \Add0~2 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~3 (
	.dataa(!mem_76_0),
	.datab(!mem_75_0),
	.datac(!mem_74_0),
	.datad(!last_packet_beat2),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add0~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~3 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~3 .lut_mask = 64'h009500FF00950000;
defparam \burst_uncompress_byte_counter~3 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[4] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[4]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[4] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[4] .power_up = "low";

cyclonev_lcell_comb \last_packet_beat~3 (
	.dataa(!\burst_uncompress_byte_counter[6]~q ),
	.datab(!\burst_uncompress_byte_counter[5]~q ),
	.datac(!\burst_uncompress_byte_counter[4]~q ),
	.datad(!\burst_uncompress_byte_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_packet_beat~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~3 .extended_lut = "off";
defparam \last_packet_beat~3 .lut_mask = 64'h8000800080008000;
defparam \last_packet_beat~3 .shared_arith = "off";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!mem_77_0),
	.datab(!mem_76_0),
	.datac(!mem_75_0),
	.datad(!mem_74_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h8000800080008000;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~6 (
	.dataa(!mem_78_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat2),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~6 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~6 .lut_mask = 64'h0000000C0A0A000C;
defparam \burst_uncompress_byte_counter~6 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[7] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[7]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[7] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[7] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[2]~q ),
	.datac(!\last_packet_beat~3_combout ),
	.datad(!\burst_uncompress_byte_counter[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~0 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~0 .lut_mask = 64'h5155515551555155;
defparam \burst_uncompress_byte_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!mem_77_0),
	.datab(!mem_76_0),
	.datac(!mem_75_0),
	.datad(!mem_74_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~2 (
	.dataa(!last_packet_beat2),
	.datab(!\burst_uncompress_byte_counter~0_combout ),
	.datac(!\Add0~1_combout ),
	.datad(!\Add1~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~2 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~2 .lut_mask = 64'h5410541054105410;
defparam \burst_uncompress_byte_counter~2 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[5] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[5]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[5] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[5] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h8000800080008000;
defparam \Add0~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~1 (
	.dataa(!mem_78_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat2),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~1 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~1 .lut_mask = 64'h0505030C0A0A030C;
defparam \burst_uncompress_byte_counter~1 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[6] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[6]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[6] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[6] .power_up = "low";

endmodule

module spw_babasu_altera_merlin_slave_agent_11 (
	h2f_RREADY_0,
	waitrequest_reset_override,
	stateST_COMP_TRANS,
	mem_used_1,
	in_data_reg_69,
	in_narrow_reg,
	wait_latency_counter_1,
	wait_latency_counter_0,
	cp_ready,
	cp_ready1,
	empty,
	mem_66_0,
	mem_used_0,
	last_packet_beat,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	last_packet_beat1,
	altera_reset_synchronizer_int_chain_out,
	last_packet_beat2,
	cp_ready2,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_RREADY_0;
input 	waitrequest_reset_override;
input 	stateST_COMP_TRANS;
input 	mem_used_1;
input 	in_data_reg_69;
input 	in_narrow_reg;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
output 	cp_ready;
output 	cp_ready1;
input 	empty;
input 	mem_66_0;
input 	mem_used_0;
output 	last_packet_beat;
input 	mem_78_0;
input 	mem_77_0;
input 	mem_76_0;
input 	mem_75_0;
input 	mem_74_0;
output 	last_packet_beat1;
input 	altera_reset_synchronizer_int_chain_out;
output 	last_packet_beat2;
output 	cp_ready2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



spw_babasu_altera_merlin_burst_uncompressor_11 uncompressor(
	.h2f_RREADY_0(h2f_RREADY_0),
	.empty(empty),
	.mem_66_0(mem_66_0),
	.mem_used_0(mem_used_0),
	.last_packet_beat(last_packet_beat),
	.mem_78_0(mem_78_0),
	.mem_77_0(mem_77_0),
	.mem_76_0(mem_76_0),
	.mem_75_0(mem_75_0),
	.mem_74_0(mem_74_0),
	.last_packet_beat1(last_packet_beat1),
	.reset(altera_reset_synchronizer_int_chain_out),
	.last_packet_beat2(last_packet_beat2),
	.clk(clk_clk));

cyclonev_lcell_comb \cp_ready~0 (
	.dataa(!waitrequest_reset_override),
	.datab(!in_data_reg_69),
	.datac(!stateST_COMP_TRANS),
	.datad(!in_narrow_reg),
	.datae(!wait_latency_counter_1),
	.dataf(!wait_latency_counter_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~0 .extended_lut = "off";
defparam \cp_ready~0 .lut_mask = 64'hCCC0CCC0DDD5CCC0;
defparam \cp_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~1 (
	.dataa(!mem_used_1),
	.datab(!cp_ready),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~1 .extended_lut = "off";
defparam \cp_ready~1 .lut_mask = 64'h2222222222222222;
defparam \cp_ready~1 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~2 (
	.dataa(!waitrequest_reset_override),
	.datab(!in_data_reg_69),
	.datac(!in_narrow_reg),
	.datad(!wait_latency_counter_1),
	.datae(!wait_latency_counter_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready2),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~2 .extended_lut = "off";
defparam \cp_ready~2 .lut_mask = 64'hC0C0D5C0C0C0D5C0;
defparam \cp_ready~2 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_burst_uncompressor_11 (
	h2f_RREADY_0,
	empty,
	mem_66_0,
	mem_used_0,
	last_packet_beat,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	last_packet_beat1,
	reset,
	last_packet_beat2,
	clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_RREADY_0;
input 	empty;
input 	mem_66_0;
input 	mem_used_0;
output 	last_packet_beat;
input 	mem_78_0;
input 	mem_77_0;
input 	mem_76_0;
input 	mem_75_0;
input 	mem_74_0;
output 	last_packet_beat1;
input 	reset;
output 	last_packet_beat2;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always0~0_combout ;
wire \burst_uncompress_busy~q ;
wire \burst_uncompress_byte_counter~5_combout ;
wire \burst_uncompress_byte_counter[2]~q ;
wire \burst_uncompress_byte_counter~4_combout ;
wire \burst_uncompress_byte_counter[3]~q ;
wire \Add0~2_combout ;
wire \burst_uncompress_byte_counter~3_combout ;
wire \burst_uncompress_byte_counter[4]~q ;
wire \last_packet_beat~3_combout ;
wire \Add1~0_combout ;
wire \burst_uncompress_byte_counter~6_combout ;
wire \burst_uncompress_byte_counter[7]~q ;
wire \burst_uncompress_byte_counter~0_combout ;
wire \Add0~1_combout ;
wire \Add1~1_combout ;
wire \burst_uncompress_byte_counter~2_combout ;
wire \burst_uncompress_byte_counter[5]~q ;
wire \Add0~0_combout ;
wire \burst_uncompress_byte_counter~1_combout ;
wire \burst_uncompress_byte_counter[6]~q ;


cyclonev_lcell_comb \last_packet_beat~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!\burst_uncompress_byte_counter[5]~q ),
	.datad(!\burst_uncompress_byte_counter[4]~q ),
	.datae(!\burst_uncompress_byte_counter[3]~q ),
	.dataf(!\burst_uncompress_byte_counter[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~0 .extended_lut = "off";
defparam \last_packet_beat~0 .lut_mask = 64'h0000000040000000;
defparam \last_packet_beat~0 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~1 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_78_0),
	.datac(!mem_77_0),
	.datad(!mem_76_0),
	.datae(!mem_75_0),
	.dataf(!mem_74_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat1),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~1 .extended_lut = "off";
defparam \last_packet_beat~1 .lut_mask = 64'h0000000080000000;
defparam \last_packet_beat~1 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~2 (
	.dataa(!empty),
	.datab(!mem_66_0),
	.datac(!mem_used_0),
	.datad(!last_packet_beat),
	.datae(!last_packet_beat1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat2),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~2 .extended_lut = "off";
defparam \last_packet_beat~2 .lut_mask = 64'h3331313133313131;
defparam \last_packet_beat~2 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!h2f_RREADY_0),
	.datab(!empty),
	.datac(!mem_used_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'h0404040404040404;
defparam \always0~0 .shared_arith = "off";

dffeas burst_uncompress_busy(
	.clk(clk),
	.d(last_packet_beat2),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_busy~q ),
	.prn(vcc));
defparam burst_uncompress_busy.is_wysiwyg = "true";
defparam burst_uncompress_busy.power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~5 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_74_0),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(!last_packet_beat2),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~5 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~5 .lut_mask = 64'h00C800FA00C800FA;
defparam \burst_uncompress_byte_counter~5 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[2] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[2]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[2] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[2] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~4 (
	.dataa(!mem_75_0),
	.datab(!mem_74_0),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(!last_packet_beat2),
	.dataf(!\burst_uncompress_byte_counter~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~4 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~4 .lut_mask = 64'h000099990000F00F;
defparam \burst_uncompress_byte_counter~4 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[3] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[3]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[3] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[3] .power_up = "low";

cyclonev_lcell_comb \Add0~2 (
	.dataa(!\burst_uncompress_byte_counter[4]~q ),
	.datab(!\burst_uncompress_byte_counter[3]~q ),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~2 .extended_lut = "off";
defparam \Add0~2 .lut_mask = 64'h6A6A6A6A6A6A6A6A;
defparam \Add0~2 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~3 (
	.dataa(!mem_76_0),
	.datab(!mem_75_0),
	.datac(!mem_74_0),
	.datad(!last_packet_beat2),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add0~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~3 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~3 .lut_mask = 64'h009500FF00950000;
defparam \burst_uncompress_byte_counter~3 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[4] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[4]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[4] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[4] .power_up = "low";

cyclonev_lcell_comb \last_packet_beat~3 (
	.dataa(!\burst_uncompress_byte_counter[6]~q ),
	.datab(!\burst_uncompress_byte_counter[5]~q ),
	.datac(!\burst_uncompress_byte_counter[4]~q ),
	.datad(!\burst_uncompress_byte_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_packet_beat~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~3 .extended_lut = "off";
defparam \last_packet_beat~3 .lut_mask = 64'h8000800080008000;
defparam \last_packet_beat~3 .shared_arith = "off";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!mem_77_0),
	.datab(!mem_76_0),
	.datac(!mem_75_0),
	.datad(!mem_74_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h8000800080008000;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~6 (
	.dataa(!mem_78_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat2),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~6 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~6 .lut_mask = 64'h0000000C0A0A000C;
defparam \burst_uncompress_byte_counter~6 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[7] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[7]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[7] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[7] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[2]~q ),
	.datac(!\last_packet_beat~3_combout ),
	.datad(!\burst_uncompress_byte_counter[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~0 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~0 .lut_mask = 64'h5155515551555155;
defparam \burst_uncompress_byte_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!mem_77_0),
	.datab(!mem_76_0),
	.datac(!mem_75_0),
	.datad(!mem_74_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~2 (
	.dataa(!last_packet_beat2),
	.datab(!\burst_uncompress_byte_counter~0_combout ),
	.datac(!\Add0~1_combout ),
	.datad(!\Add1~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~2 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~2 .lut_mask = 64'h5410541054105410;
defparam \burst_uncompress_byte_counter~2 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[5] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[5]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[5] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[5] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h8000800080008000;
defparam \Add0~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~1 (
	.dataa(!mem_78_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat2),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~1 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~1 .lut_mask = 64'h0505030C0A0A030C;
defparam \burst_uncompress_byte_counter~1 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[6] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[6]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[6] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[6] .power_up = "low";

endmodule

module spw_babasu_altera_merlin_slave_agent_12 (
	waitrequest_reset_override,
	stateST_COMP_TRANS,
	out_valid_reg,
	mem_used_1,
	in_narrow_reg,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	WideOr0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	in_data_reg_68,
	cp_ready,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_129_0,
	mem_used_01,
	mem_66_0,
	comb,
	last_packet_beat,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	last_packet_beat1,
	altera_reset_synchronizer_int_chain_out,
	m0_write1,
	nxt_out_eop,
	cp_ready1,
	last_packet_beat2,
	read,
	cp_ready2,
	in_data_reg_69,
	rf_source_valid,
	rp_valid1,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	waitrequest_reset_override;
input 	stateST_COMP_TRANS;
input 	out_valid_reg;
input 	mem_used_1;
input 	in_narrow_reg;
input 	in_byteen_reg_3;
input 	in_byteen_reg_2;
input 	in_byteen_reg_1;
input 	in_byteen_reg_0;
output 	WideOr0;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	in_data_reg_68;
output 	cp_ready;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	mem_129_0;
input 	mem_used_01;
input 	mem_66_0;
output 	comb;
output 	last_packet_beat;
input 	mem_78_0;
input 	mem_77_0;
input 	mem_76_0;
input 	mem_75_0;
input 	mem_74_0;
output 	last_packet_beat1;
input 	altera_reset_synchronizer_int_chain_out;
output 	m0_write1;
input 	nxt_out_eop;
output 	cp_ready1;
output 	last_packet_beat2;
input 	read;
output 	cp_ready2;
input 	in_data_reg_69;
output 	rf_source_valid;
output 	rp_valid1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \local_write~combout ;
wire \cp_ready~1_combout ;
wire \cp_ready~2_combout ;


spw_babasu_altera_merlin_burst_uncompressor_12 uncompressor(
	.mem_66_0(mem_66_0),
	.comb(comb),
	.last_packet_beat(last_packet_beat),
	.mem_78_0(mem_78_0),
	.mem_77_0(mem_77_0),
	.mem_76_0(mem_76_0),
	.mem_75_0(mem_75_0),
	.mem_74_0(mem_74_0),
	.last_packet_beat1(last_packet_beat1),
	.reset(altera_reset_synchronizer_int_chain_out),
	.last_packet_beat2(last_packet_beat2),
	.read(read),
	.clk(clk_clk));

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!in_narrow_reg),
	.datac(!in_byteen_reg_3),
	.datad(!in_byteen_reg_2),
	.datae(!in_byteen_reg_1),
	.dataf(!in_byteen_reg_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h1FFFFFFFFFFFFFFF;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~0 (
	.dataa(!waitrequest_reset_override),
	.datab(!mem_used_1),
	.datac(!WideOr0),
	.datad(!wait_latency_counter_1),
	.datae(!wait_latency_counter_0),
	.dataf(!\local_write~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~0 .extended_lut = "off";
defparam \cp_ready~0 .lut_mask = 64'hC0C0C4C0C4C0C0C0;
defparam \cp_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \comb~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_129_0),
	.datad(!mem_used_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(comb),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~0 .extended_lut = "off";
defparam \comb~0 .lut_mask = 64'h007F007F007F007F;
defparam \comb~0 .shared_arith = "off";

cyclonev_lcell_comb m0_write(
	.dataa(!mem_used_1),
	.datab(!WideOr0),
	.datac(!\local_write~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write1),
	.sumout(),
	.cout(),
	.shareout());
defparam m0_write.extended_lut = "off";
defparam m0_write.lut_mask = 64'h0202020202020202;
defparam m0_write.shared_arith = "off";

cyclonev_lcell_comb \cp_ready~3 (
	.dataa(!mem_used_1),
	.datab(!in_narrow_reg),
	.datac(!\cp_ready~1_combout ),
	.datad(!\cp_ready~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~3 .extended_lut = "off";
defparam \cp_ready~3 .lut_mask = 64'h08AA08AA08AA08AA;
defparam \cp_ready~3 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~4 (
	.dataa(!waitrequest_reset_override),
	.datab(!mem_used_1),
	.datac(!WideOr0),
	.datad(!wait_latency_counter_1),
	.datae(!wait_latency_counter_0),
	.dataf(!\local_write~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready2),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~4 .extended_lut = "off";
defparam \cp_ready~4 .lut_mask = 64'h0000550004005100;
defparam \cp_ready~4 .shared_arith = "off";

cyclonev_lcell_comb \rf_source_valid~0 (
	.dataa(!in_data_reg_68),
	.datab(!out_valid_reg),
	.datac(!nxt_out_eop),
	.datad(!in_data_reg_69),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rf_source_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_source_valid~0 .extended_lut = "off";
defparam \rf_source_valid~0 .lut_mask = 64'h0133013301330133;
defparam \rf_source_valid~0 .shared_arith = "off";

cyclonev_lcell_comb rp_valid(
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_129_0),
	.datad(!mem_used_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rp_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam rp_valid.extended_lut = "off";
defparam rp_valid.lut_mask = 64'h8880888088808880;
defparam rp_valid.shared_arith = "off";

cyclonev_lcell_comb local_write(
	.dataa(!in_data_reg_68),
	.datab(!out_valid_reg),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\local_write~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam local_write.extended_lut = "off";
defparam local_write.lut_mask = 64'h1111111111111111;
defparam local_write.shared_arith = "off";

cyclonev_lcell_comb \cp_ready~1 (
	.dataa(!in_byteen_reg_3),
	.datab(!in_byteen_reg_2),
	.datac(!in_byteen_reg_1),
	.datad(!in_byteen_reg_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cp_ready~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~1 .extended_lut = "off";
defparam \cp_ready~1 .lut_mask = 64'h8000800080008000;
defparam \cp_ready~1 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~2 (
	.dataa(!waitrequest_reset_override),
	.datab(!wait_latency_counter_1),
	.datac(!wait_latency_counter_0),
	.datad(!\local_write~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cp_ready~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~2 .extended_lut = "off";
defparam \cp_ready~2 .lut_mask = 64'h0440044004400440;
defparam \cp_ready~2 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_burst_uncompressor_12 (
	mem_66_0,
	comb,
	last_packet_beat,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	last_packet_beat1,
	reset,
	last_packet_beat2,
	read,
	clk)/* synthesis synthesis_greybox=0 */;
input 	mem_66_0;
input 	comb;
output 	last_packet_beat;
input 	mem_78_0;
input 	mem_77_0;
input 	mem_76_0;
input 	mem_75_0;
input 	mem_74_0;
output 	last_packet_beat1;
input 	reset;
output 	last_packet_beat2;
input 	read;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \burst_uncompress_busy~q ;
wire \burst_uncompress_byte_counter~5_combout ;
wire \burst_uncompress_byte_counter[2]~q ;
wire \burst_uncompress_byte_counter~4_combout ;
wire \burst_uncompress_byte_counter[3]~q ;
wire \Add0~2_combout ;
wire \burst_uncompress_byte_counter~3_combout ;
wire \burst_uncompress_byte_counter[4]~q ;
wire \last_packet_beat~3_combout ;
wire \Add1~0_combout ;
wire \burst_uncompress_byte_counter~6_combout ;
wire \burst_uncompress_byte_counter[7]~q ;
wire \burst_uncompress_byte_counter~0_combout ;
wire \Add0~1_combout ;
wire \Add1~1_combout ;
wire \burst_uncompress_byte_counter~2_combout ;
wire \burst_uncompress_byte_counter[5]~q ;
wire \Add0~0_combout ;
wire \burst_uncompress_byte_counter~1_combout ;
wire \burst_uncompress_byte_counter[6]~q ;


cyclonev_lcell_comb \last_packet_beat~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!\burst_uncompress_byte_counter[5]~q ),
	.datad(!\burst_uncompress_byte_counter[4]~q ),
	.datae(!\burst_uncompress_byte_counter[3]~q ),
	.dataf(!\burst_uncompress_byte_counter[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~0 .extended_lut = "off";
defparam \last_packet_beat~0 .lut_mask = 64'h0000000040000000;
defparam \last_packet_beat~0 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~1 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_78_0),
	.datac(!mem_77_0),
	.datad(!mem_76_0),
	.datae(!mem_75_0),
	.dataf(!mem_74_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat1),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~1 .extended_lut = "off";
defparam \last_packet_beat~1 .lut_mask = 64'h0000000080000000;
defparam \last_packet_beat~1 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~2 (
	.dataa(!comb),
	.datab(!mem_66_0),
	.datac(!last_packet_beat),
	.datad(!last_packet_beat1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat2),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~2 .extended_lut = "off";
defparam \last_packet_beat~2 .lut_mask = 64'h3222322232223222;
defparam \last_packet_beat~2 .shared_arith = "off";

dffeas burst_uncompress_busy(
	.clk(clk),
	.d(last_packet_beat2),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_busy~q ),
	.prn(vcc));
defparam burst_uncompress_busy.is_wysiwyg = "true";
defparam burst_uncompress_busy.power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~5 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_74_0),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(!last_packet_beat2),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~5 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~5 .lut_mask = 64'h00C800FA00C800FA;
defparam \burst_uncompress_byte_counter~5 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[2] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[2]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[2] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[2] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~4 (
	.dataa(!mem_75_0),
	.datab(!mem_74_0),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(!last_packet_beat2),
	.dataf(!\burst_uncompress_byte_counter~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~4 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~4 .lut_mask = 64'h000099990000F00F;
defparam \burst_uncompress_byte_counter~4 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[3] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[3]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[3] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[3] .power_up = "low";

cyclonev_lcell_comb \Add0~2 (
	.dataa(!\burst_uncompress_byte_counter[4]~q ),
	.datab(!\burst_uncompress_byte_counter[3]~q ),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~2 .extended_lut = "off";
defparam \Add0~2 .lut_mask = 64'h6A6A6A6A6A6A6A6A;
defparam \Add0~2 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~3 (
	.dataa(!mem_76_0),
	.datab(!mem_75_0),
	.datac(!mem_74_0),
	.datad(!last_packet_beat2),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add0~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~3 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~3 .lut_mask = 64'h009500FF00950000;
defparam \burst_uncompress_byte_counter~3 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[4] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[4]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[4] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[4] .power_up = "low";

cyclonev_lcell_comb \last_packet_beat~3 (
	.dataa(!\burst_uncompress_byte_counter[6]~q ),
	.datab(!\burst_uncompress_byte_counter[5]~q ),
	.datac(!\burst_uncompress_byte_counter[4]~q ),
	.datad(!\burst_uncompress_byte_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_packet_beat~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~3 .extended_lut = "off";
defparam \last_packet_beat~3 .lut_mask = 64'h8000800080008000;
defparam \last_packet_beat~3 .shared_arith = "off";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!mem_77_0),
	.datab(!mem_76_0),
	.datac(!mem_75_0),
	.datad(!mem_74_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h8000800080008000;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~6 (
	.dataa(!mem_78_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat2),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~6 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~6 .lut_mask = 64'h0000000C0A0A000C;
defparam \burst_uncompress_byte_counter~6 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[7] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[7]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[7] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[7] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[2]~q ),
	.datac(!\last_packet_beat~3_combout ),
	.datad(!\burst_uncompress_byte_counter[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~0 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~0 .lut_mask = 64'h5155515551555155;
defparam \burst_uncompress_byte_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!mem_77_0),
	.datab(!mem_76_0),
	.datac(!mem_75_0),
	.datad(!mem_74_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~2 (
	.dataa(!last_packet_beat2),
	.datab(!\burst_uncompress_byte_counter~0_combout ),
	.datac(!\Add0~1_combout ),
	.datad(!\Add1~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~2 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~2 .lut_mask = 64'h5410541054105410;
defparam \burst_uncompress_byte_counter~2 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[5] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[5]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[5] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[5] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h8000800080008000;
defparam \Add0~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~1 (
	.dataa(!mem_78_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat2),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~1 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~1 .lut_mask = 64'h0505030C0A0A030C;
defparam \burst_uncompress_byte_counter~1 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[6] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[6]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[6] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[6] .power_up = "low";

endmodule

module spw_babasu_altera_merlin_slave_agent_13 (
	h2f_RREADY_0,
	waitrequest_reset_override,
	stateST_COMP_TRANS,
	mem_used_1,
	in_data_reg_69,
	in_narrow_reg,
	wait_latency_counter_1,
	wait_latency_counter_0,
	cp_ready,
	cp_ready1,
	empty,
	mem_66_0,
	mem_used_0,
	last_packet_beat,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	last_packet_beat1,
	altera_reset_synchronizer_int_chain_out,
	last_packet_beat2,
	cp_ready2,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_RREADY_0;
input 	waitrequest_reset_override;
input 	stateST_COMP_TRANS;
input 	mem_used_1;
input 	in_data_reg_69;
input 	in_narrow_reg;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
output 	cp_ready;
output 	cp_ready1;
input 	empty;
input 	mem_66_0;
input 	mem_used_0;
output 	last_packet_beat;
input 	mem_78_0;
input 	mem_77_0;
input 	mem_76_0;
input 	mem_75_0;
input 	mem_74_0;
output 	last_packet_beat1;
input 	altera_reset_synchronizer_int_chain_out;
output 	last_packet_beat2;
output 	cp_ready2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



spw_babasu_altera_merlin_burst_uncompressor_13 uncompressor(
	.h2f_RREADY_0(h2f_RREADY_0),
	.empty(empty),
	.mem_66_0(mem_66_0),
	.mem_used_0(mem_used_0),
	.last_packet_beat(last_packet_beat),
	.mem_78_0(mem_78_0),
	.mem_77_0(mem_77_0),
	.mem_76_0(mem_76_0),
	.mem_75_0(mem_75_0),
	.mem_74_0(mem_74_0),
	.last_packet_beat1(last_packet_beat1),
	.reset(altera_reset_synchronizer_int_chain_out),
	.last_packet_beat2(last_packet_beat2),
	.clk(clk_clk));

cyclonev_lcell_comb \cp_ready~0 (
	.dataa(!waitrequest_reset_override),
	.datab(!in_data_reg_69),
	.datac(!stateST_COMP_TRANS),
	.datad(!in_narrow_reg),
	.datae(!wait_latency_counter_1),
	.dataf(!wait_latency_counter_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~0 .extended_lut = "off";
defparam \cp_ready~0 .lut_mask = 64'hCCC0CCC0DDD5CCC0;
defparam \cp_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~1 (
	.dataa(!mem_used_1),
	.datab(!cp_ready),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~1 .extended_lut = "off";
defparam \cp_ready~1 .lut_mask = 64'h2222222222222222;
defparam \cp_ready~1 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~2 (
	.dataa(!waitrequest_reset_override),
	.datab(!in_data_reg_69),
	.datac(!in_narrow_reg),
	.datad(!wait_latency_counter_1),
	.datae(!wait_latency_counter_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready2),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~2 .extended_lut = "off";
defparam \cp_ready~2 .lut_mask = 64'hC0C0D5C0C0C0D5C0;
defparam \cp_ready~2 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_burst_uncompressor_13 (
	h2f_RREADY_0,
	empty,
	mem_66_0,
	mem_used_0,
	last_packet_beat,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	last_packet_beat1,
	reset,
	last_packet_beat2,
	clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_RREADY_0;
input 	empty;
input 	mem_66_0;
input 	mem_used_0;
output 	last_packet_beat;
input 	mem_78_0;
input 	mem_77_0;
input 	mem_76_0;
input 	mem_75_0;
input 	mem_74_0;
output 	last_packet_beat1;
input 	reset;
output 	last_packet_beat2;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always0~0_combout ;
wire \burst_uncompress_busy~q ;
wire \burst_uncompress_byte_counter~5_combout ;
wire \burst_uncompress_byte_counter[2]~q ;
wire \burst_uncompress_byte_counter~4_combout ;
wire \burst_uncompress_byte_counter[3]~q ;
wire \Add0~2_combout ;
wire \burst_uncompress_byte_counter~3_combout ;
wire \burst_uncompress_byte_counter[4]~q ;
wire \last_packet_beat~3_combout ;
wire \Add1~0_combout ;
wire \burst_uncompress_byte_counter~6_combout ;
wire \burst_uncompress_byte_counter[7]~q ;
wire \burst_uncompress_byte_counter~0_combout ;
wire \Add0~1_combout ;
wire \Add1~1_combout ;
wire \burst_uncompress_byte_counter~2_combout ;
wire \burst_uncompress_byte_counter[5]~q ;
wire \Add0~0_combout ;
wire \burst_uncompress_byte_counter~1_combout ;
wire \burst_uncompress_byte_counter[6]~q ;


cyclonev_lcell_comb \last_packet_beat~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!\burst_uncompress_byte_counter[5]~q ),
	.datad(!\burst_uncompress_byte_counter[4]~q ),
	.datae(!\burst_uncompress_byte_counter[3]~q ),
	.dataf(!\burst_uncompress_byte_counter[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~0 .extended_lut = "off";
defparam \last_packet_beat~0 .lut_mask = 64'h0000000040000000;
defparam \last_packet_beat~0 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~1 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_78_0),
	.datac(!mem_77_0),
	.datad(!mem_76_0),
	.datae(!mem_75_0),
	.dataf(!mem_74_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat1),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~1 .extended_lut = "off";
defparam \last_packet_beat~1 .lut_mask = 64'h0000000080000000;
defparam \last_packet_beat~1 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~2 (
	.dataa(!empty),
	.datab(!mem_66_0),
	.datac(!mem_used_0),
	.datad(!last_packet_beat),
	.datae(!last_packet_beat1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat2),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~2 .extended_lut = "off";
defparam \last_packet_beat~2 .lut_mask = 64'h3331313133313131;
defparam \last_packet_beat~2 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!h2f_RREADY_0),
	.datab(!empty),
	.datac(!mem_used_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'h0404040404040404;
defparam \always0~0 .shared_arith = "off";

dffeas burst_uncompress_busy(
	.clk(clk),
	.d(last_packet_beat2),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_busy~q ),
	.prn(vcc));
defparam burst_uncompress_busy.is_wysiwyg = "true";
defparam burst_uncompress_busy.power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~5 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_74_0),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(!last_packet_beat2),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~5 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~5 .lut_mask = 64'h00C800FA00C800FA;
defparam \burst_uncompress_byte_counter~5 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[2] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[2]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[2] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[2] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~4 (
	.dataa(!mem_75_0),
	.datab(!mem_74_0),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(!last_packet_beat2),
	.dataf(!\burst_uncompress_byte_counter~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~4 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~4 .lut_mask = 64'h000099990000F00F;
defparam \burst_uncompress_byte_counter~4 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[3] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[3]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[3] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[3] .power_up = "low";

cyclonev_lcell_comb \Add0~2 (
	.dataa(!\burst_uncompress_byte_counter[4]~q ),
	.datab(!\burst_uncompress_byte_counter[3]~q ),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~2 .extended_lut = "off";
defparam \Add0~2 .lut_mask = 64'h6A6A6A6A6A6A6A6A;
defparam \Add0~2 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~3 (
	.dataa(!mem_76_0),
	.datab(!mem_75_0),
	.datac(!mem_74_0),
	.datad(!last_packet_beat2),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add0~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~3 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~3 .lut_mask = 64'h009500FF00950000;
defparam \burst_uncompress_byte_counter~3 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[4] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[4]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[4] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[4] .power_up = "low";

cyclonev_lcell_comb \last_packet_beat~3 (
	.dataa(!\burst_uncompress_byte_counter[6]~q ),
	.datab(!\burst_uncompress_byte_counter[5]~q ),
	.datac(!\burst_uncompress_byte_counter[4]~q ),
	.datad(!\burst_uncompress_byte_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_packet_beat~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~3 .extended_lut = "off";
defparam \last_packet_beat~3 .lut_mask = 64'h8000800080008000;
defparam \last_packet_beat~3 .shared_arith = "off";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!mem_77_0),
	.datab(!mem_76_0),
	.datac(!mem_75_0),
	.datad(!mem_74_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h8000800080008000;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~6 (
	.dataa(!mem_78_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat2),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~6 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~6 .lut_mask = 64'h0000000C0A0A000C;
defparam \burst_uncompress_byte_counter~6 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[7] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[7]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[7] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[7] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[2]~q ),
	.datac(!\last_packet_beat~3_combout ),
	.datad(!\burst_uncompress_byte_counter[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~0 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~0 .lut_mask = 64'h5155515551555155;
defparam \burst_uncompress_byte_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!mem_77_0),
	.datab(!mem_76_0),
	.datac(!mem_75_0),
	.datad(!mem_74_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~2 (
	.dataa(!last_packet_beat2),
	.datab(!\burst_uncompress_byte_counter~0_combout ),
	.datac(!\Add0~1_combout ),
	.datad(!\Add1~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~2 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~2 .lut_mask = 64'h5410541054105410;
defparam \burst_uncompress_byte_counter~2 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[5] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[5]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[5] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[5] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h8000800080008000;
defparam \Add0~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~1 (
	.dataa(!mem_78_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat2),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~1 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~1 .lut_mask = 64'h0505030C0A0A030C;
defparam \burst_uncompress_byte_counter~1 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[6] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[6]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[6] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[6] .power_up = "low";

endmodule

module spw_babasu_altera_merlin_slave_agent_14 (
	waitrequest_reset_override,
	stateST_COMP_TRANS,
	out_valid_reg,
	mem_used_1,
	in_narrow_reg,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	WideOr0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	in_data_reg_68,
	cp_ready,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_129_0,
	mem_used_01,
	mem_66_0,
	comb,
	last_packet_beat,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	last_packet_beat1,
	altera_reset_synchronizer_int_chain_out,
	m0_write1,
	nxt_out_eop,
	cp_ready1,
	last_packet_beat2,
	WideOr01,
	read,
	cp_ready2,
	in_data_reg_69,
	rf_source_valid,
	rf_sink_ready,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	waitrequest_reset_override;
input 	stateST_COMP_TRANS;
input 	out_valid_reg;
input 	mem_used_1;
input 	in_narrow_reg;
input 	in_byteen_reg_3;
input 	in_byteen_reg_2;
input 	in_byteen_reg_1;
input 	in_byteen_reg_0;
output 	WideOr0;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	in_data_reg_68;
output 	cp_ready;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	mem_129_0;
input 	mem_used_01;
input 	mem_66_0;
output 	comb;
output 	last_packet_beat;
input 	mem_78_0;
input 	mem_77_0;
input 	mem_76_0;
input 	mem_75_0;
input 	mem_74_0;
output 	last_packet_beat1;
input 	altera_reset_synchronizer_int_chain_out;
output 	m0_write1;
input 	nxt_out_eop;
output 	cp_ready1;
output 	last_packet_beat2;
input 	WideOr01;
input 	read;
output 	cp_ready2;
input 	in_data_reg_69;
output 	rf_source_valid;
output 	rf_sink_ready;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \local_write~combout ;
wire \cp_ready~1_combout ;
wire \cp_ready~2_combout ;


spw_babasu_altera_merlin_burst_uncompressor_14 uncompressor(
	.mem_66_0(mem_66_0),
	.comb(comb),
	.last_packet_beat(last_packet_beat),
	.mem_78_0(mem_78_0),
	.mem_77_0(mem_77_0),
	.mem_76_0(mem_76_0),
	.mem_75_0(mem_75_0),
	.mem_74_0(mem_74_0),
	.last_packet_beat1(last_packet_beat1),
	.reset(altera_reset_synchronizer_int_chain_out),
	.last_packet_beat2(last_packet_beat2),
	.WideOr0(WideOr01),
	.read(read),
	.sink_ready(rf_sink_ready),
	.clk(clk_clk));

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!in_narrow_reg),
	.datac(!in_byteen_reg_3),
	.datad(!in_byteen_reg_2),
	.datae(!in_byteen_reg_1),
	.dataf(!in_byteen_reg_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h1FFFFFFFFFFFFFFF;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~0 (
	.dataa(!waitrequest_reset_override),
	.datab(!mem_used_1),
	.datac(!WideOr0),
	.datad(!wait_latency_counter_1),
	.datae(!wait_latency_counter_0),
	.dataf(!\local_write~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~0 .extended_lut = "off";
defparam \cp_ready~0 .lut_mask = 64'hC0C0C4C0C4C0C0C0;
defparam \cp_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \comb~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_129_0),
	.datad(!mem_used_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(comb),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~0 .extended_lut = "off";
defparam \comb~0 .lut_mask = 64'h007F007F007F007F;
defparam \comb~0 .shared_arith = "off";

cyclonev_lcell_comb m0_write(
	.dataa(!mem_used_1),
	.datab(!WideOr0),
	.datac(!\local_write~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write1),
	.sumout(),
	.cout(),
	.shareout());
defparam m0_write.extended_lut = "off";
defparam m0_write.lut_mask = 64'h0202020202020202;
defparam m0_write.shared_arith = "off";

cyclonev_lcell_comb \cp_ready~3 (
	.dataa(!mem_used_1),
	.datab(!in_narrow_reg),
	.datac(!\cp_ready~1_combout ),
	.datad(!\cp_ready~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~3 .extended_lut = "off";
defparam \cp_ready~3 .lut_mask = 64'h08AA08AA08AA08AA;
defparam \cp_ready~3 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~4 (
	.dataa(!waitrequest_reset_override),
	.datab(!mem_used_1),
	.datac(!WideOr0),
	.datad(!wait_latency_counter_1),
	.datae(!wait_latency_counter_0),
	.dataf(!\local_write~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready2),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~4 .extended_lut = "off";
defparam \cp_ready~4 .lut_mask = 64'h0000550004005100;
defparam \cp_ready~4 .shared_arith = "off";

cyclonev_lcell_comb \rf_source_valid~0 (
	.dataa(!in_data_reg_68),
	.datab(!out_valid_reg),
	.datac(!nxt_out_eop),
	.datad(!in_data_reg_69),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rf_source_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_source_valid~0 .extended_lut = "off";
defparam \rf_source_valid~0 .lut_mask = 64'h0133013301330133;
defparam \rf_source_valid~0 .shared_arith = "off";

cyclonev_lcell_comb local_write(
	.dataa(!in_data_reg_68),
	.datab(!out_valid_reg),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\local_write~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam local_write.extended_lut = "off";
defparam local_write.lut_mask = 64'h1111111111111111;
defparam local_write.shared_arith = "off";

cyclonev_lcell_comb \cp_ready~1 (
	.dataa(!in_byteen_reg_3),
	.datab(!in_byteen_reg_2),
	.datac(!in_byteen_reg_1),
	.datad(!in_byteen_reg_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cp_ready~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~1 .extended_lut = "off";
defparam \cp_ready~1 .lut_mask = 64'h8000800080008000;
defparam \cp_ready~1 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~2 (
	.dataa(!waitrequest_reset_override),
	.datab(!wait_latency_counter_1),
	.datac(!wait_latency_counter_0),
	.datad(!\local_write~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cp_ready~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~2 .extended_lut = "off";
defparam \cp_ready~2 .lut_mask = 64'h0440044004400440;
defparam \cp_ready~2 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_burst_uncompressor_14 (
	mem_66_0,
	comb,
	last_packet_beat,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	last_packet_beat1,
	reset,
	last_packet_beat2,
	WideOr0,
	read,
	sink_ready,
	clk)/* synthesis synthesis_greybox=0 */;
input 	mem_66_0;
input 	comb;
output 	last_packet_beat;
input 	mem_78_0;
input 	mem_77_0;
input 	mem_76_0;
input 	mem_75_0;
input 	mem_74_0;
output 	last_packet_beat1;
input 	reset;
output 	last_packet_beat2;
input 	WideOr0;
input 	read;
output 	sink_ready;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \burst_uncompress_busy~q ;
wire \burst_uncompress_byte_counter~5_combout ;
wire \burst_uncompress_byte_counter[2]~q ;
wire \burst_uncompress_byte_counter~4_combout ;
wire \burst_uncompress_byte_counter[3]~q ;
wire \Add0~2_combout ;
wire \burst_uncompress_byte_counter~3_combout ;
wire \burst_uncompress_byte_counter[4]~q ;
wire \last_packet_beat~3_combout ;
wire \Add1~0_combout ;
wire \burst_uncompress_byte_counter~6_combout ;
wire \burst_uncompress_byte_counter[7]~q ;
wire \burst_uncompress_byte_counter~0_combout ;
wire \Add0~1_combout ;
wire \Add1~1_combout ;
wire \burst_uncompress_byte_counter~2_combout ;
wire \burst_uncompress_byte_counter[5]~q ;
wire \Add0~0_combout ;
wire \burst_uncompress_byte_counter~1_combout ;
wire \burst_uncompress_byte_counter[6]~q ;


cyclonev_lcell_comb \last_packet_beat~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!\burst_uncompress_byte_counter[5]~q ),
	.datad(!\burst_uncompress_byte_counter[4]~q ),
	.datae(!\burst_uncompress_byte_counter[3]~q ),
	.dataf(!\burst_uncompress_byte_counter[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~0 .extended_lut = "off";
defparam \last_packet_beat~0 .lut_mask = 64'h0000000040000000;
defparam \last_packet_beat~0 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~1 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_78_0),
	.datac(!mem_77_0),
	.datad(!mem_76_0),
	.datae(!mem_75_0),
	.dataf(!mem_74_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat1),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~1 .extended_lut = "off";
defparam \last_packet_beat~1 .lut_mask = 64'h0000000080000000;
defparam \last_packet_beat~1 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~2 (
	.dataa(!comb),
	.datab(!mem_66_0),
	.datac(!last_packet_beat),
	.datad(!last_packet_beat1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat2),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~2 .extended_lut = "off";
defparam \last_packet_beat~2 .lut_mask = 64'h3222322232223222;
defparam \last_packet_beat~2 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!comb),
	.datad(!last_packet_beat2),
	.datae(!WideOr0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~0 .extended_lut = "off";
defparam \sink_ready~0 .lut_mask = 64'h00000F0000000F00;
defparam \sink_ready~0 .shared_arith = "off";

dffeas burst_uncompress_busy(
	.clk(clk),
	.d(last_packet_beat2),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_busy~q ),
	.prn(vcc));
defparam burst_uncompress_busy.is_wysiwyg = "true";
defparam burst_uncompress_busy.power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~5 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_74_0),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(!last_packet_beat2),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~5 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~5 .lut_mask = 64'h00C800FA00C800FA;
defparam \burst_uncompress_byte_counter~5 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[2] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[2]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[2] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[2] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~4 (
	.dataa(!mem_75_0),
	.datab(!mem_74_0),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(!last_packet_beat2),
	.dataf(!\burst_uncompress_byte_counter~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~4 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~4 .lut_mask = 64'h000099990000F00F;
defparam \burst_uncompress_byte_counter~4 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[3] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[3]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[3] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[3] .power_up = "low";

cyclonev_lcell_comb \Add0~2 (
	.dataa(!\burst_uncompress_byte_counter[4]~q ),
	.datab(!\burst_uncompress_byte_counter[3]~q ),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~2 .extended_lut = "off";
defparam \Add0~2 .lut_mask = 64'h6A6A6A6A6A6A6A6A;
defparam \Add0~2 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~3 (
	.dataa(!mem_76_0),
	.datab(!mem_75_0),
	.datac(!mem_74_0),
	.datad(!last_packet_beat2),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add0~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~3 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~3 .lut_mask = 64'h009500FF00950000;
defparam \burst_uncompress_byte_counter~3 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[4] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[4]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[4] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[4] .power_up = "low";

cyclonev_lcell_comb \last_packet_beat~3 (
	.dataa(!\burst_uncompress_byte_counter[6]~q ),
	.datab(!\burst_uncompress_byte_counter[5]~q ),
	.datac(!\burst_uncompress_byte_counter[4]~q ),
	.datad(!\burst_uncompress_byte_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_packet_beat~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~3 .extended_lut = "off";
defparam \last_packet_beat~3 .lut_mask = 64'h8000800080008000;
defparam \last_packet_beat~3 .shared_arith = "off";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!mem_77_0),
	.datab(!mem_76_0),
	.datac(!mem_75_0),
	.datad(!mem_74_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h8000800080008000;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~6 (
	.dataa(!mem_78_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat2),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~6 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~6 .lut_mask = 64'h0000000C0A0A000C;
defparam \burst_uncompress_byte_counter~6 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[7] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[7]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[7] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[7] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[2]~q ),
	.datac(!\last_packet_beat~3_combout ),
	.datad(!\burst_uncompress_byte_counter[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~0 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~0 .lut_mask = 64'h5155515551555155;
defparam \burst_uncompress_byte_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!mem_77_0),
	.datab(!mem_76_0),
	.datac(!mem_75_0),
	.datad(!mem_74_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~2 (
	.dataa(!last_packet_beat2),
	.datab(!\burst_uncompress_byte_counter~0_combout ),
	.datac(!\Add0~1_combout ),
	.datad(!\Add1~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~2 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~2 .lut_mask = 64'h5410541054105410;
defparam \burst_uncompress_byte_counter~2 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[5] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[5]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[5] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[5] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h8000800080008000;
defparam \Add0~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~1 (
	.dataa(!mem_78_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat2),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~1 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~1 .lut_mask = 64'h0505030C0A0A030C;
defparam \burst_uncompress_byte_counter~1 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[6] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[6]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[6] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[6] .power_up = "low";

endmodule

module spw_babasu_altera_merlin_slave_agent_15 (
	h2f_RREADY_0,
	waitrequest_reset_override,
	in_data_reg_69,
	stateST_COMP_TRANS,
	in_narrow_reg,
	wait_latency_counter_1,
	wait_latency_counter_0,
	cp_ready,
	empty,
	mem_66_0,
	mem_used_0,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	last_packet_beat,
	altera_reset_synchronizer_int_chain_out,
	cp_ready1,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_RREADY_0;
input 	waitrequest_reset_override;
input 	in_data_reg_69;
input 	stateST_COMP_TRANS;
input 	in_narrow_reg;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
output 	cp_ready;
input 	empty;
input 	mem_66_0;
input 	mem_used_0;
input 	mem_78_0;
input 	mem_77_0;
input 	mem_76_0;
input 	mem_75_0;
input 	mem_74_0;
output 	last_packet_beat;
input 	altera_reset_synchronizer_int_chain_out;
output 	cp_ready1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



spw_babasu_altera_merlin_burst_uncompressor_15 uncompressor(
	.h2f_RREADY_0(h2f_RREADY_0),
	.empty(empty),
	.mem_66_0(mem_66_0),
	.mem_used_0(mem_used_0),
	.mem_78_0(mem_78_0),
	.mem_77_0(mem_77_0),
	.mem_76_0(mem_76_0),
	.mem_75_0(mem_75_0),
	.mem_74_0(mem_74_0),
	.last_packet_beat(last_packet_beat),
	.reset(altera_reset_synchronizer_int_chain_out),
	.clk(clk_clk));

cyclonev_lcell_comb \cp_ready~0 (
	.dataa(!waitrequest_reset_override),
	.datab(!in_data_reg_69),
	.datac(!stateST_COMP_TRANS),
	.datad(!in_narrow_reg),
	.datae(!wait_latency_counter_1),
	.dataf(!wait_latency_counter_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~0 .extended_lut = "off";
defparam \cp_ready~0 .lut_mask = 64'hCCC0CCC0DDD5CCC0;
defparam \cp_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~1 (
	.dataa(!waitrequest_reset_override),
	.datab(!in_data_reg_69),
	.datac(!in_narrow_reg),
	.datad(!wait_latency_counter_1),
	.datae(!wait_latency_counter_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~1 .extended_lut = "off";
defparam \cp_ready~1 .lut_mask = 64'hC0C0D5C0C0C0D5C0;
defparam \cp_ready~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_burst_uncompressor_15 (
	h2f_RREADY_0,
	empty,
	mem_66_0,
	mem_used_0,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	last_packet_beat,
	reset,
	clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_RREADY_0;
input 	empty;
input 	mem_66_0;
input 	mem_used_0;
input 	mem_78_0;
input 	mem_77_0;
input 	mem_76_0;
input 	mem_75_0;
input 	mem_74_0;
output 	last_packet_beat;
input 	reset;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always0~0_combout ;
wire \burst_uncompress_busy~q ;
wire \burst_uncompress_byte_counter~5_combout ;
wire \burst_uncompress_byte_counter[3]~q ;
wire \Add0~2_combout ;
wire \burst_uncompress_byte_counter~4_combout ;
wire \burst_uncompress_byte_counter[4]~q ;
wire \Add0~1_combout ;
wire \Add1~1_combout ;
wire \burst_uncompress_byte_counter~3_combout ;
wire \burst_uncompress_byte_counter[5]~q ;
wire \Add0~0_combout ;
wire \Add1~0_combout ;
wire \burst_uncompress_byte_counter~2_combout ;
wire \burst_uncompress_byte_counter[6]~q ;
wire \last_packet_beat~1_combout ;
wire \burst_uncompress_byte_counter~6_combout ;
wire \burst_uncompress_byte_counter[7]~q ;
wire \burst_uncompress_byte_counter~0_combout ;
wire \burst_uncompress_byte_counter~1_combout ;
wire \burst_uncompress_byte_counter[2]~q ;
wire \last_packet_beat~0_combout ;
wire \last_packet_beat~2_combout ;


cyclonev_lcell_comb \last_packet_beat~3 (
	.dataa(!empty),
	.datab(!mem_66_0),
	.datac(!mem_used_0),
	.datad(!\last_packet_beat~0_combout ),
	.datae(!\last_packet_beat~1_combout ),
	.dataf(!\last_packet_beat~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~3 .extended_lut = "off";
defparam \last_packet_beat~3 .lut_mask = 64'h3333333131313131;
defparam \last_packet_beat~3 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!h2f_RREADY_0),
	.datab(!empty),
	.datac(!mem_used_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'h0404040404040404;
defparam \always0~0 .shared_arith = "off";

dffeas burst_uncompress_busy(
	.clk(clk),
	.d(last_packet_beat),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_busy~q ),
	.prn(vcc));
defparam burst_uncompress_busy.is_wysiwyg = "true";
defparam burst_uncompress_busy.power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~5 (
	.dataa(!mem_75_0),
	.datab(!mem_74_0),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(!last_packet_beat),
	.dataf(!\burst_uncompress_byte_counter~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~5 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~5 .lut_mask = 64'h000099990000F00F;
defparam \burst_uncompress_byte_counter~5 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[3] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[3]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[3] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[3] .power_up = "low";

cyclonev_lcell_comb \Add0~2 (
	.dataa(!\burst_uncompress_byte_counter[4]~q ),
	.datab(!\burst_uncompress_byte_counter[3]~q ),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~2 .extended_lut = "off";
defparam \Add0~2 .lut_mask = 64'h6A6A6A6A6A6A6A6A;
defparam \Add0~2 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~4 (
	.dataa(!mem_76_0),
	.datab(!mem_75_0),
	.datac(!mem_74_0),
	.datad(!last_packet_beat),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add0~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~4 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~4 .lut_mask = 64'h009500FF00950000;
defparam \burst_uncompress_byte_counter~4 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[4] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[4]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[4] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[4] .power_up = "low";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!mem_77_0),
	.datab(!mem_76_0),
	.datac(!mem_75_0),
	.datad(!mem_74_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~3 (
	.dataa(!last_packet_beat),
	.datab(!\burst_uncompress_byte_counter~0_combout ),
	.datac(!\Add0~1_combout ),
	.datad(!\Add1~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~3 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~3 .lut_mask = 64'h5410541054105410;
defparam \burst_uncompress_byte_counter~3 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[5] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[5]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[5] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[5] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h8000800080008000;
defparam \Add0~0 .shared_arith = "off";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!mem_77_0),
	.datab(!mem_76_0),
	.datac(!mem_75_0),
	.datad(!mem_74_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h8000800080008000;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~2 (
	.dataa(!mem_78_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~2 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~2 .lut_mask = 64'h0505030C0A0A030C;
defparam \burst_uncompress_byte_counter~2 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[6] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[6]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[6] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[6] .power_up = "low";

cyclonev_lcell_comb \last_packet_beat~1 (
	.dataa(!\burst_uncompress_byte_counter[6]~q ),
	.datab(!\burst_uncompress_byte_counter[5]~q ),
	.datac(!\burst_uncompress_byte_counter[4]~q ),
	.datad(!\burst_uncompress_byte_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_packet_beat~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~1 .extended_lut = "off";
defparam \last_packet_beat~1 .lut_mask = 64'h8000800080008000;
defparam \last_packet_beat~1 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~6 (
	.dataa(!mem_78_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~6 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~6 .lut_mask = 64'h0000000C0A0A000C;
defparam \burst_uncompress_byte_counter~6 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[7] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[7]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[7] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[7] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[2]~q ),
	.datac(!\last_packet_beat~1_combout ),
	.datad(!\burst_uncompress_byte_counter[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~0 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~0 .lut_mask = 64'h5155515551555155;
defparam \burst_uncompress_byte_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~1 (
	.dataa(!mem_74_0),
	.datab(!\last_packet_beat~0_combout ),
	.datac(!last_packet_beat),
	.datad(!\burst_uncompress_byte_counter~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~1 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~1 .lut_mask = 64'h080C080C080C080C;
defparam \burst_uncompress_byte_counter~1 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[2] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[2]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[2] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[2] .power_up = "low";

cyclonev_lcell_comb \last_packet_beat~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_packet_beat~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~0 .extended_lut = "off";
defparam \last_packet_beat~0 .lut_mask = 64'h1111111111111111;
defparam \last_packet_beat~0 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~2 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_78_0),
	.datac(!mem_77_0),
	.datad(!mem_76_0),
	.datae(!mem_75_0),
	.dataf(!mem_74_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_packet_beat~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~2 .extended_lut = "off";
defparam \last_packet_beat~2 .lut_mask = 64'h0000000080000000;
defparam \last_packet_beat~2 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_slave_agent_16 (
	waitrequest_reset_override,
	stateST_COMP_TRANS,
	out_valid_reg,
	mem_used_1,
	in_narrow_reg,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	WideOr0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	in_data_reg_68,
	cp_ready,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_129_0,
	mem_used_01,
	mem_66_0,
	comb,
	last_packet_beat,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	last_packet_beat1,
	altera_reset_synchronizer_int_chain_out,
	m0_write1,
	nxt_out_eop,
	cp_ready1,
	last_packet_beat2,
	WideOr01,
	read,
	cp_ready2,
	in_data_reg_69,
	rf_source_valid,
	rf_sink_ready,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	waitrequest_reset_override;
input 	stateST_COMP_TRANS;
input 	out_valid_reg;
input 	mem_used_1;
input 	in_narrow_reg;
input 	in_byteen_reg_3;
input 	in_byteen_reg_2;
input 	in_byteen_reg_1;
input 	in_byteen_reg_0;
output 	WideOr0;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	in_data_reg_68;
output 	cp_ready;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	mem_129_0;
input 	mem_used_01;
input 	mem_66_0;
output 	comb;
output 	last_packet_beat;
input 	mem_78_0;
input 	mem_77_0;
input 	mem_76_0;
input 	mem_75_0;
input 	mem_74_0;
output 	last_packet_beat1;
input 	altera_reset_synchronizer_int_chain_out;
output 	m0_write1;
input 	nxt_out_eop;
output 	cp_ready1;
output 	last_packet_beat2;
input 	WideOr01;
input 	read;
output 	cp_ready2;
input 	in_data_reg_69;
output 	rf_source_valid;
output 	rf_sink_ready;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \local_write~combout ;
wire \cp_ready~1_combout ;
wire \cp_ready~2_combout ;


spw_babasu_altera_merlin_burst_uncompressor_16 uncompressor(
	.mem_66_0(mem_66_0),
	.comb(comb),
	.last_packet_beat(last_packet_beat),
	.mem_78_0(mem_78_0),
	.mem_77_0(mem_77_0),
	.mem_76_0(mem_76_0),
	.mem_75_0(mem_75_0),
	.mem_74_0(mem_74_0),
	.last_packet_beat1(last_packet_beat1),
	.reset(altera_reset_synchronizer_int_chain_out),
	.last_packet_beat2(last_packet_beat2),
	.WideOr0(WideOr01),
	.read(read),
	.sink_ready(rf_sink_ready),
	.clk(clk_clk));

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!in_narrow_reg),
	.datac(!in_byteen_reg_3),
	.datad(!in_byteen_reg_2),
	.datae(!in_byteen_reg_1),
	.dataf(!in_byteen_reg_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h1FFFFFFFFFFFFFFF;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~0 (
	.dataa(!waitrequest_reset_override),
	.datab(!mem_used_1),
	.datac(!WideOr0),
	.datad(!wait_latency_counter_1),
	.datae(!wait_latency_counter_0),
	.dataf(!\local_write~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~0 .extended_lut = "off";
defparam \cp_ready~0 .lut_mask = 64'hC0C0C4C0C4C0C0C0;
defparam \cp_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \comb~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_129_0),
	.datad(!mem_used_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(comb),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~0 .extended_lut = "off";
defparam \comb~0 .lut_mask = 64'h007F007F007F007F;
defparam \comb~0 .shared_arith = "off";

cyclonev_lcell_comb m0_write(
	.dataa(!mem_used_1),
	.datab(!WideOr0),
	.datac(!\local_write~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write1),
	.sumout(),
	.cout(),
	.shareout());
defparam m0_write.extended_lut = "off";
defparam m0_write.lut_mask = 64'h0202020202020202;
defparam m0_write.shared_arith = "off";

cyclonev_lcell_comb \cp_ready~3 (
	.dataa(!mem_used_1),
	.datab(!in_narrow_reg),
	.datac(!\cp_ready~1_combout ),
	.datad(!\cp_ready~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~3 .extended_lut = "off";
defparam \cp_ready~3 .lut_mask = 64'h08AA08AA08AA08AA;
defparam \cp_ready~3 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~4 (
	.dataa(!waitrequest_reset_override),
	.datab(!mem_used_1),
	.datac(!WideOr0),
	.datad(!wait_latency_counter_1),
	.datae(!wait_latency_counter_0),
	.dataf(!\local_write~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready2),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~4 .extended_lut = "off";
defparam \cp_ready~4 .lut_mask = 64'h0000550004005100;
defparam \cp_ready~4 .shared_arith = "off";

cyclonev_lcell_comb \rf_source_valid~0 (
	.dataa(!in_data_reg_68),
	.datab(!out_valid_reg),
	.datac(!nxt_out_eop),
	.datad(!in_data_reg_69),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rf_source_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_source_valid~0 .extended_lut = "off";
defparam \rf_source_valid~0 .lut_mask = 64'h0133013301330133;
defparam \rf_source_valid~0 .shared_arith = "off";

cyclonev_lcell_comb local_write(
	.dataa(!in_data_reg_68),
	.datab(!out_valid_reg),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\local_write~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam local_write.extended_lut = "off";
defparam local_write.lut_mask = 64'h1111111111111111;
defparam local_write.shared_arith = "off";

cyclonev_lcell_comb \cp_ready~1 (
	.dataa(!in_byteen_reg_3),
	.datab(!in_byteen_reg_2),
	.datac(!in_byteen_reg_1),
	.datad(!in_byteen_reg_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cp_ready~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~1 .extended_lut = "off";
defparam \cp_ready~1 .lut_mask = 64'h8000800080008000;
defparam \cp_ready~1 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~2 (
	.dataa(!waitrequest_reset_override),
	.datab(!wait_latency_counter_1),
	.datac(!wait_latency_counter_0),
	.datad(!\local_write~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cp_ready~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~2 .extended_lut = "off";
defparam \cp_ready~2 .lut_mask = 64'h0440044004400440;
defparam \cp_ready~2 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_burst_uncompressor_16 (
	mem_66_0,
	comb,
	last_packet_beat,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	last_packet_beat1,
	reset,
	last_packet_beat2,
	WideOr0,
	read,
	sink_ready,
	clk)/* synthesis synthesis_greybox=0 */;
input 	mem_66_0;
input 	comb;
output 	last_packet_beat;
input 	mem_78_0;
input 	mem_77_0;
input 	mem_76_0;
input 	mem_75_0;
input 	mem_74_0;
output 	last_packet_beat1;
input 	reset;
output 	last_packet_beat2;
input 	WideOr0;
input 	read;
output 	sink_ready;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \burst_uncompress_busy~q ;
wire \burst_uncompress_byte_counter~5_combout ;
wire \burst_uncompress_byte_counter[2]~q ;
wire \burst_uncompress_byte_counter~4_combout ;
wire \burst_uncompress_byte_counter[3]~q ;
wire \Add0~2_combout ;
wire \burst_uncompress_byte_counter~3_combout ;
wire \burst_uncompress_byte_counter[4]~q ;
wire \last_packet_beat~3_combout ;
wire \Add1~0_combout ;
wire \burst_uncompress_byte_counter~6_combout ;
wire \burst_uncompress_byte_counter[7]~q ;
wire \burst_uncompress_byte_counter~0_combout ;
wire \Add0~1_combout ;
wire \Add1~1_combout ;
wire \burst_uncompress_byte_counter~2_combout ;
wire \burst_uncompress_byte_counter[5]~q ;
wire \Add0~0_combout ;
wire \burst_uncompress_byte_counter~1_combout ;
wire \burst_uncompress_byte_counter[6]~q ;


cyclonev_lcell_comb \last_packet_beat~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!\burst_uncompress_byte_counter[5]~q ),
	.datad(!\burst_uncompress_byte_counter[4]~q ),
	.datae(!\burst_uncompress_byte_counter[3]~q ),
	.dataf(!\burst_uncompress_byte_counter[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~0 .extended_lut = "off";
defparam \last_packet_beat~0 .lut_mask = 64'h0000000040000000;
defparam \last_packet_beat~0 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~1 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_78_0),
	.datac(!mem_77_0),
	.datad(!mem_76_0),
	.datae(!mem_75_0),
	.dataf(!mem_74_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat1),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~1 .extended_lut = "off";
defparam \last_packet_beat~1 .lut_mask = 64'h0000000080000000;
defparam \last_packet_beat~1 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~2 (
	.dataa(!comb),
	.datab(!mem_66_0),
	.datac(!last_packet_beat),
	.datad(!last_packet_beat1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat2),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~2 .extended_lut = "off";
defparam \last_packet_beat~2 .lut_mask = 64'h3222322232223222;
defparam \last_packet_beat~2 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!comb),
	.datad(!last_packet_beat2),
	.datae(!WideOr0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~0 .extended_lut = "off";
defparam \sink_ready~0 .lut_mask = 64'h00000F0000000F00;
defparam \sink_ready~0 .shared_arith = "off";

dffeas burst_uncompress_busy(
	.clk(clk),
	.d(last_packet_beat2),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_busy~q ),
	.prn(vcc));
defparam burst_uncompress_busy.is_wysiwyg = "true";
defparam burst_uncompress_busy.power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~5 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_74_0),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(!last_packet_beat2),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~5 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~5 .lut_mask = 64'h00C800FA00C800FA;
defparam \burst_uncompress_byte_counter~5 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[2] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[2]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[2] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[2] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~4 (
	.dataa(!mem_75_0),
	.datab(!mem_74_0),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(!last_packet_beat2),
	.dataf(!\burst_uncompress_byte_counter~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~4 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~4 .lut_mask = 64'h000099990000F00F;
defparam \burst_uncompress_byte_counter~4 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[3] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[3]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[3] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[3] .power_up = "low";

cyclonev_lcell_comb \Add0~2 (
	.dataa(!\burst_uncompress_byte_counter[4]~q ),
	.datab(!\burst_uncompress_byte_counter[3]~q ),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~2 .extended_lut = "off";
defparam \Add0~2 .lut_mask = 64'h6A6A6A6A6A6A6A6A;
defparam \Add0~2 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~3 (
	.dataa(!mem_76_0),
	.datab(!mem_75_0),
	.datac(!mem_74_0),
	.datad(!last_packet_beat2),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add0~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~3 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~3 .lut_mask = 64'h009500FF00950000;
defparam \burst_uncompress_byte_counter~3 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[4] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[4]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[4] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[4] .power_up = "low";

cyclonev_lcell_comb \last_packet_beat~3 (
	.dataa(!\burst_uncompress_byte_counter[6]~q ),
	.datab(!\burst_uncompress_byte_counter[5]~q ),
	.datac(!\burst_uncompress_byte_counter[4]~q ),
	.datad(!\burst_uncompress_byte_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_packet_beat~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~3 .extended_lut = "off";
defparam \last_packet_beat~3 .lut_mask = 64'h8000800080008000;
defparam \last_packet_beat~3 .shared_arith = "off";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!mem_77_0),
	.datab(!mem_76_0),
	.datac(!mem_75_0),
	.datad(!mem_74_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h8000800080008000;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~6 (
	.dataa(!mem_78_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat2),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~6 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~6 .lut_mask = 64'h0000000C0A0A000C;
defparam \burst_uncompress_byte_counter~6 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[7] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[7]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[7] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[7] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[2]~q ),
	.datac(!\last_packet_beat~3_combout ),
	.datad(!\burst_uncompress_byte_counter[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~0 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~0 .lut_mask = 64'h5155515551555155;
defparam \burst_uncompress_byte_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!mem_77_0),
	.datab(!mem_76_0),
	.datac(!mem_75_0),
	.datad(!mem_74_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~2 (
	.dataa(!last_packet_beat2),
	.datab(!\burst_uncompress_byte_counter~0_combout ),
	.datac(!\Add0~1_combout ),
	.datad(!\Add1~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~2 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~2 .lut_mask = 64'h5410541054105410;
defparam \burst_uncompress_byte_counter~2 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[5] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[5]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[5] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[5] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h8000800080008000;
defparam \Add0~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~1 (
	.dataa(!mem_78_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat2),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~1 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~1 .lut_mask = 64'h0505030C0A0A030C;
defparam \burst_uncompress_byte_counter~1 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[6] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[6]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[6] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[6] .power_up = "low";

endmodule

module spw_babasu_altera_merlin_slave_translator (
	waitrequest_reset_override1,
	out_valid_reg,
	mem_used_1,
	WideOr0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	read_latency_shift_reg_0,
	av_readdata_pre_0,
	m0_write,
	reset,
	cp_ready,
	in_data_reg_69,
	av_readdata,
	clk)/* synthesis synthesis_greybox=0 */;
output 	waitrequest_reset_override1;
input 	out_valid_reg;
input 	mem_used_1;
input 	WideOr0;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
output 	read_latency_shift_reg_0;
output 	av_readdata_pre_0;
input 	m0_write;
input 	reset;
input 	cp_ready;
input 	in_data_reg_69;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~0_combout ;
wire \wait_latency_counter[0]~0_combout ;
wire \wait_latency_counter~1_combout ;
wire \wait_latency_counter~2_combout ;
wire \read_latency_shift_reg~1_combout ;


dffeas waitrequest_reset_override(
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(waitrequest_reset_override1),
	.prn(vcc));
defparam waitrequest_reset_override.is_wysiwyg = "true";
defparam waitrequest_reset_override.power_up = "low";

dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!mem_used_1),
	.datab(!WideOr0),
	.datac(!out_valid_reg),
	.datad(!in_data_reg_69),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'h0002000200020002;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter[0]~0 (
	.dataa(!waitrequest_reset_override1),
	.datab(!wait_latency_counter_1),
	.datac(!wait_latency_counter_0),
	.datad(!m0_write),
	.datae(!\read_latency_shift_reg~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter[0]~0 .extended_lut = "off";
defparam \wait_latency_counter[0]~0 .lut_mask = 64'h0015511500155115;
defparam \wait_latency_counter[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!\wait_latency_counter[0]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'h0606060606060606;
defparam \wait_latency_counter~1 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~2 (
	.dataa(!wait_latency_counter_0),
	.datab(!\wait_latency_counter[0]~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~2 .extended_lut = "off";
defparam \wait_latency_counter~2 .lut_mask = 64'h2222222222222222;
defparam \wait_latency_counter~2 .shared_arith = "off";

cyclonev_lcell_comb \read_latency_shift_reg~1 (
	.dataa(!cp_ready),
	.datab(!\read_latency_shift_reg~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~1 .extended_lut = "off";
defparam \read_latency_shift_reg~1 .lut_mask = 64'h1111111111111111;
defparam \read_latency_shift_reg~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_slave_translator_1 (
	wait_latency_counter_1,
	wait_latency_counter_0,
	read_latency_shift_reg_0,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	reset,
	write,
	write1,
	av_readdata,
	clk)/* synthesis synthesis_greybox=0 */;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
output 	read_latency_shift_reg_0;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
input 	reset;
input 	write;
input 	write1;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter~0_combout ;
wire \wait_latency_counter~1_combout ;


dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(write1),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

cyclonev_lcell_comb \wait_latency_counter~0 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!write),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~0 .extended_lut = "off";
defparam \wait_latency_counter~0 .lut_mask = 64'h0404040404040404;
defparam \wait_latency_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(gnd),
	.datab(!wait_latency_counter_0),
	.datac(!write),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'h0C0C0C0C0C0C0C0C;
defparam \wait_latency_counter~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_slave_translator_2 (
	waitrequest_reset_override,
	out_valid_reg,
	mem_used_1,
	WideOr0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	read_latency_shift_reg_0,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata_pre_7,
	av_readdata_pre_8,
	reset,
	m0_write,
	cp_ready,
	in_data_reg_69,
	av_readdata,
	clk)/* synthesis synthesis_greybox=0 */;
input 	waitrequest_reset_override;
input 	out_valid_reg;
input 	mem_used_1;
input 	WideOr0;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
output 	read_latency_shift_reg_0;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
output 	av_readdata_pre_6;
output 	av_readdata_pre_7;
output 	av_readdata_pre_8;
input 	reset;
input 	m0_write;
input 	cp_ready;
input 	in_data_reg_69;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~0_combout ;
wire \wait_latency_counter[1]~0_combout ;
wire \wait_latency_counter~1_combout ;
wire \wait_latency_counter~2_combout ;
wire \read_latency_shift_reg~1_combout ;


dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!mem_used_1),
	.datab(!WideOr0),
	.datac(!out_valid_reg),
	.datad(!in_data_reg_69),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'h0002000200020002;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter[1]~0 (
	.dataa(!waitrequest_reset_override),
	.datab(!wait_latency_counter_1),
	.datac(!wait_latency_counter_0),
	.datad(!m0_write),
	.datae(!\read_latency_shift_reg~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter[1]~0 .extended_lut = "off";
defparam \wait_latency_counter[1]~0 .lut_mask = 64'h0015511500155115;
defparam \wait_latency_counter[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!\wait_latency_counter[1]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'h0606060606060606;
defparam \wait_latency_counter~1 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~2 (
	.dataa(!wait_latency_counter_0),
	.datab(!\wait_latency_counter[1]~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~2 .extended_lut = "off";
defparam \wait_latency_counter~2 .lut_mask = 64'h2222222222222222;
defparam \wait_latency_counter~2 .shared_arith = "off";

cyclonev_lcell_comb \read_latency_shift_reg~1 (
	.dataa(!cp_ready),
	.datab(!\read_latency_shift_reg~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~1 .extended_lut = "off";
defparam \read_latency_shift_reg~1 .lut_mask = 64'h1111111111111111;
defparam \read_latency_shift_reg~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_slave_translator_3 (
	wait_latency_counter_1,
	wait_latency_counter_0,
	read_latency_shift_reg_0,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata_pre_7,
	av_readdata_pre_8,
	reset,
	write,
	write1,
	av_readdata,
	clk)/* synthesis synthesis_greybox=0 */;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
output 	read_latency_shift_reg_0;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
output 	av_readdata_pre_6;
output 	av_readdata_pre_7;
output 	av_readdata_pre_8;
input 	reset;
input 	write;
input 	write1;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter~0_combout ;
wire \wait_latency_counter~1_combout ;


dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(write1),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

cyclonev_lcell_comb \wait_latency_counter~0 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!write),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~0 .extended_lut = "off";
defparam \wait_latency_counter~0 .lut_mask = 64'h0404040404040404;
defparam \wait_latency_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(gnd),
	.datab(!wait_latency_counter_0),
	.datac(!write),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'h0C0C0C0C0C0C0C0C;
defparam \wait_latency_counter~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_slave_translator_4 (
	wait_latency_counter_1,
	wait_latency_counter_0,
	read_latency_shift_reg_0,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata_pre_7,
	av_readdata_pre_8,
	av_readdata_pre_9,
	av_readdata_pre_10,
	reset,
	write,
	write1,
	av_readdata,
	clk)/* synthesis synthesis_greybox=0 */;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
output 	read_latency_shift_reg_0;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
output 	av_readdata_pre_6;
output 	av_readdata_pre_7;
output 	av_readdata_pre_8;
output 	av_readdata_pre_9;
output 	av_readdata_pre_10;
input 	reset;
input 	write;
input 	write1;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter~0_combout ;
wire \wait_latency_counter~1_combout ;


dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(write1),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

dffeas \av_readdata_pre[9] (
	.clk(clk),
	.d(av_readdata[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_9),
	.prn(vcc));
defparam \av_readdata_pre[9] .is_wysiwyg = "true";
defparam \av_readdata_pre[9] .power_up = "low";

dffeas \av_readdata_pre[10] (
	.clk(clk),
	.d(av_readdata[10]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_10),
	.prn(vcc));
defparam \av_readdata_pre[10] .is_wysiwyg = "true";
defparam \av_readdata_pre[10] .power_up = "low";

cyclonev_lcell_comb \wait_latency_counter~0 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!write),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~0 .extended_lut = "off";
defparam \wait_latency_counter~0 .lut_mask = 64'h0404040404040404;
defparam \wait_latency_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(gnd),
	.datab(!wait_latency_counter_0),
	.datac(!write),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'h0C0C0C0C0C0C0C0C;
defparam \wait_latency_counter~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_slave_translator_5 (
	waitrequest_reset_override,
	out_valid_reg,
	mem_used_1,
	WideOr0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	read_latency_shift_reg_0,
	av_readdata_pre_0,
	reset,
	m0_write,
	cp_ready,
	in_data_reg_69,
	av_readdata,
	clk)/* synthesis synthesis_greybox=0 */;
input 	waitrequest_reset_override;
input 	out_valid_reg;
input 	mem_used_1;
input 	WideOr0;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
output 	read_latency_shift_reg_0;
output 	av_readdata_pre_0;
input 	reset;
input 	m0_write;
input 	cp_ready;
input 	in_data_reg_69;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~0_combout ;
wire \wait_latency_counter[1]~0_combout ;
wire \wait_latency_counter~1_combout ;
wire \wait_latency_counter~2_combout ;
wire \read_latency_shift_reg~1_combout ;


dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!mem_used_1),
	.datab(!WideOr0),
	.datac(!out_valid_reg),
	.datad(!in_data_reg_69),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'h0002000200020002;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter[1]~0 (
	.dataa(!waitrequest_reset_override),
	.datab(!wait_latency_counter_1),
	.datac(!wait_latency_counter_0),
	.datad(!m0_write),
	.datae(!\read_latency_shift_reg~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter[1]~0 .extended_lut = "off";
defparam \wait_latency_counter[1]~0 .lut_mask = 64'h0015511500155115;
defparam \wait_latency_counter[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!\wait_latency_counter[1]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'h0606060606060606;
defparam \wait_latency_counter~1 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~2 (
	.dataa(!wait_latency_counter_0),
	.datab(!\wait_latency_counter[1]~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~2 .extended_lut = "off";
defparam \wait_latency_counter~2 .lut_mask = 64'h2222222222222222;
defparam \wait_latency_counter~2 .shared_arith = "off";

cyclonev_lcell_comb \read_latency_shift_reg~1 (
	.dataa(!cp_ready),
	.datab(!\read_latency_shift_reg~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~1 .extended_lut = "off";
defparam \read_latency_shift_reg~1 .lut_mask = 64'h1111111111111111;
defparam \read_latency_shift_reg~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_slave_translator_6 (
	waitrequest_reset_override,
	out_valid_reg,
	mem_used_1,
	WideOr0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	read_latency_shift_reg_0,
	av_readdata_pre_0,
	reset,
	m0_write,
	cp_ready,
	in_data_reg_69,
	av_readdata,
	clk)/* synthesis synthesis_greybox=0 */;
input 	waitrequest_reset_override;
input 	out_valid_reg;
input 	mem_used_1;
input 	WideOr0;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
output 	read_latency_shift_reg_0;
output 	av_readdata_pre_0;
input 	reset;
input 	m0_write;
input 	cp_ready;
input 	in_data_reg_69;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~0_combout ;
wire \wait_latency_counter[1]~0_combout ;
wire \wait_latency_counter~1_combout ;
wire \wait_latency_counter~2_combout ;
wire \read_latency_shift_reg~1_combout ;


dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!mem_used_1),
	.datab(!WideOr0),
	.datac(!out_valid_reg),
	.datad(!in_data_reg_69),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'h0002000200020002;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter[1]~0 (
	.dataa(!waitrequest_reset_override),
	.datab(!wait_latency_counter_1),
	.datac(!wait_latency_counter_0),
	.datad(!m0_write),
	.datae(!\read_latency_shift_reg~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter[1]~0 .extended_lut = "off";
defparam \wait_latency_counter[1]~0 .lut_mask = 64'h0015511500155115;
defparam \wait_latency_counter[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!\wait_latency_counter[1]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'h0606060606060606;
defparam \wait_latency_counter~1 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~2 (
	.dataa(!wait_latency_counter_0),
	.datab(!\wait_latency_counter[1]~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~2 .extended_lut = "off";
defparam \wait_latency_counter~2 .lut_mask = 64'h2222222222222222;
defparam \wait_latency_counter~2 .shared_arith = "off";

cyclonev_lcell_comb \read_latency_shift_reg~1 (
	.dataa(!cp_ready),
	.datab(!\read_latency_shift_reg~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~1 .extended_lut = "off";
defparam \read_latency_shift_reg~1 .lut_mask = 64'h1111111111111111;
defparam \read_latency_shift_reg~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_slave_translator_7 (
	waitrequest_reset_override,
	out_valid_reg,
	mem_used_1,
	WideOr0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	read_latency_shift_reg_0,
	av_readdata_pre_0,
	reset,
	m0_write,
	cp_ready,
	in_data_reg_69,
	av_readdata,
	clk)/* synthesis synthesis_greybox=0 */;
input 	waitrequest_reset_override;
input 	out_valid_reg;
input 	mem_used_1;
input 	WideOr0;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
output 	read_latency_shift_reg_0;
output 	av_readdata_pre_0;
input 	reset;
input 	m0_write;
input 	cp_ready;
input 	in_data_reg_69;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~0_combout ;
wire \wait_latency_counter[1]~0_combout ;
wire \wait_latency_counter~1_combout ;
wire \wait_latency_counter~2_combout ;
wire \read_latency_shift_reg~1_combout ;


dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!mem_used_1),
	.datab(!WideOr0),
	.datac(!out_valid_reg),
	.datad(!in_data_reg_69),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'h0002000200020002;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter[1]~0 (
	.dataa(!waitrequest_reset_override),
	.datab(!wait_latency_counter_1),
	.datac(!wait_latency_counter_0),
	.datad(!m0_write),
	.datae(!\read_latency_shift_reg~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter[1]~0 .extended_lut = "off";
defparam \wait_latency_counter[1]~0 .lut_mask = 64'h0015511500155115;
defparam \wait_latency_counter[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!\wait_latency_counter[1]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'h0606060606060606;
defparam \wait_latency_counter~1 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~2 (
	.dataa(!wait_latency_counter_0),
	.datab(!\wait_latency_counter[1]~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~2 .extended_lut = "off";
defparam \wait_latency_counter~2 .lut_mask = 64'h2222222222222222;
defparam \wait_latency_counter~2 .shared_arith = "off";

cyclonev_lcell_comb \read_latency_shift_reg~1 (
	.dataa(!cp_ready),
	.datab(!\read_latency_shift_reg~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~1 .extended_lut = "off";
defparam \read_latency_shift_reg~1 .lut_mask = 64'h1111111111111111;
defparam \read_latency_shift_reg~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_slave_translator_8 (
	wait_latency_counter_1,
	wait_latency_counter_0,
	read_latency_shift_reg_0,
	av_readdata_pre_0,
	reset,
	write,
	write1,
	av_readdata,
	clk)/* synthesis synthesis_greybox=0 */;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
output 	read_latency_shift_reg_0;
output 	av_readdata_pre_0;
input 	reset;
input 	write;
input 	write1;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter~0_combout ;
wire \wait_latency_counter~1_combout ;


dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(write1),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

cyclonev_lcell_comb \wait_latency_counter~0 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!write),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~0 .extended_lut = "off";
defparam \wait_latency_counter~0 .lut_mask = 64'h0404040404040404;
defparam \wait_latency_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(gnd),
	.datab(!wait_latency_counter_0),
	.datac(!write),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'h0C0C0C0C0C0C0C0C;
defparam \wait_latency_counter~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_slave_translator_9 (
	waitrequest_reset_override,
	out_valid_reg,
	mem_used_1,
	WideOr0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	read_latency_shift_reg_0,
	av_readdata_pre_0,
	reset,
	m0_write,
	cp_ready,
	in_data_reg_69,
	av_readdata,
	clk)/* synthesis synthesis_greybox=0 */;
input 	waitrequest_reset_override;
input 	out_valid_reg;
input 	mem_used_1;
input 	WideOr0;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
output 	read_latency_shift_reg_0;
output 	av_readdata_pre_0;
input 	reset;
input 	m0_write;
input 	cp_ready;
input 	in_data_reg_69;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~0_combout ;
wire \wait_latency_counter[0]~0_combout ;
wire \wait_latency_counter~1_combout ;
wire \wait_latency_counter~2_combout ;
wire \read_latency_shift_reg~1_combout ;


dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!mem_used_1),
	.datab(!WideOr0),
	.datac(!out_valid_reg),
	.datad(!in_data_reg_69),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'h0002000200020002;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter[0]~0 (
	.dataa(!waitrequest_reset_override),
	.datab(!wait_latency_counter_1),
	.datac(!wait_latency_counter_0),
	.datad(!m0_write),
	.datae(!\read_latency_shift_reg~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter[0]~0 .extended_lut = "off";
defparam \wait_latency_counter[0]~0 .lut_mask = 64'h0015511500155115;
defparam \wait_latency_counter[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!\wait_latency_counter[0]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'h0606060606060606;
defparam \wait_latency_counter~1 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~2 (
	.dataa(!wait_latency_counter_0),
	.datab(!\wait_latency_counter[0]~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~2 .extended_lut = "off";
defparam \wait_latency_counter~2 .lut_mask = 64'h2222222222222222;
defparam \wait_latency_counter~2 .shared_arith = "off";

cyclonev_lcell_comb \read_latency_shift_reg~1 (
	.dataa(!cp_ready),
	.datab(!\read_latency_shift_reg~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~1 .extended_lut = "off";
defparam \read_latency_shift_reg~1 .lut_mask = 64'h1111111111111111;
defparam \read_latency_shift_reg~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_slave_translator_10 (
	waitrequest_reset_override,
	out_valid_reg,
	mem_used_1,
	WideOr0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	read_latency_shift_reg_0,
	av_readdata_pre_0,
	reset,
	m0_write,
	cp_ready,
	in_data_reg_69,
	av_readdata,
	clk)/* synthesis synthesis_greybox=0 */;
input 	waitrequest_reset_override;
input 	out_valid_reg;
input 	mem_used_1;
input 	WideOr0;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
output 	read_latency_shift_reg_0;
output 	av_readdata_pre_0;
input 	reset;
input 	m0_write;
input 	cp_ready;
input 	in_data_reg_69;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~0_combout ;
wire \wait_latency_counter[0]~0_combout ;
wire \wait_latency_counter~1_combout ;
wire \wait_latency_counter~2_combout ;
wire \read_latency_shift_reg~1_combout ;


dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!mem_used_1),
	.datab(!WideOr0),
	.datac(!out_valid_reg),
	.datad(!in_data_reg_69),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'h0002000200020002;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter[0]~0 (
	.dataa(!waitrequest_reset_override),
	.datab(!wait_latency_counter_1),
	.datac(!wait_latency_counter_0),
	.datad(!m0_write),
	.datae(!\read_latency_shift_reg~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter[0]~0 .extended_lut = "off";
defparam \wait_latency_counter[0]~0 .lut_mask = 64'h0015511500155115;
defparam \wait_latency_counter[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!\wait_latency_counter[0]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'h0606060606060606;
defparam \wait_latency_counter~1 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~2 (
	.dataa(!wait_latency_counter_0),
	.datab(!\wait_latency_counter[0]~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~2 .extended_lut = "off";
defparam \wait_latency_counter~2 .lut_mask = 64'h2222222222222222;
defparam \wait_latency_counter~2 .shared_arith = "off";

cyclonev_lcell_comb \read_latency_shift_reg~1 (
	.dataa(!cp_ready),
	.datab(!\read_latency_shift_reg~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~1 .extended_lut = "off";
defparam \read_latency_shift_reg~1 .lut_mask = 64'h1111111111111111;
defparam \read_latency_shift_reg~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_slave_translator_11 (
	wait_latency_counter_1,
	wait_latency_counter_0,
	read_latency_shift_reg_0,
	av_readdata_pre_0,
	reset,
	write,
	write1,
	av_readdata,
	clk)/* synthesis synthesis_greybox=0 */;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
output 	read_latency_shift_reg_0;
output 	av_readdata_pre_0;
input 	reset;
input 	write;
input 	write1;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter~0_combout ;
wire \wait_latency_counter~1_combout ;


dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(write1),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

cyclonev_lcell_comb \wait_latency_counter~0 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!write),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~0 .extended_lut = "off";
defparam \wait_latency_counter~0 .lut_mask = 64'h0404040404040404;
defparam \wait_latency_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(gnd),
	.datab(!wait_latency_counter_0),
	.datac(!write),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'h0C0C0C0C0C0C0C0C;
defparam \wait_latency_counter~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_slave_translator_12 (
	waitrequest_reset_override,
	out_valid_reg,
	mem_used_1,
	WideOr0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	read_latency_shift_reg_0,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata_pre_7,
	reset,
	m0_write,
	cp_ready,
	in_data_reg_69,
	av_readdata,
	clk)/* synthesis synthesis_greybox=0 */;
input 	waitrequest_reset_override;
input 	out_valid_reg;
input 	mem_used_1;
input 	WideOr0;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
output 	read_latency_shift_reg_0;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
output 	av_readdata_pre_6;
output 	av_readdata_pre_7;
input 	reset;
input 	m0_write;
input 	cp_ready;
input 	in_data_reg_69;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~0_combout ;
wire \wait_latency_counter[0]~0_combout ;
wire \wait_latency_counter~1_combout ;
wire \wait_latency_counter~2_combout ;
wire \read_latency_shift_reg~1_combout ;


dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!mem_used_1),
	.datab(!WideOr0),
	.datac(!out_valid_reg),
	.datad(!in_data_reg_69),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'h0002000200020002;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter[0]~0 (
	.dataa(!waitrequest_reset_override),
	.datab(!wait_latency_counter_1),
	.datac(!wait_latency_counter_0),
	.datad(!m0_write),
	.datae(!\read_latency_shift_reg~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter[0]~0 .extended_lut = "off";
defparam \wait_latency_counter[0]~0 .lut_mask = 64'h0015511500155115;
defparam \wait_latency_counter[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!\wait_latency_counter[0]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'h0606060606060606;
defparam \wait_latency_counter~1 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~2 (
	.dataa(!wait_latency_counter_0),
	.datab(!\wait_latency_counter[0]~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~2 .extended_lut = "off";
defparam \wait_latency_counter~2 .lut_mask = 64'h2222222222222222;
defparam \wait_latency_counter~2 .shared_arith = "off";

cyclonev_lcell_comb \read_latency_shift_reg~1 (
	.dataa(!cp_ready),
	.datab(!\read_latency_shift_reg~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~1 .extended_lut = "off";
defparam \read_latency_shift_reg~1 .lut_mask = 64'h1111111111111111;
defparam \read_latency_shift_reg~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_slave_translator_13 (
	wait_latency_counter_1,
	wait_latency_counter_0,
	read_latency_shift_reg_0,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata_pre_7,
	reset,
	write,
	write1,
	av_readdata,
	clk)/* synthesis synthesis_greybox=0 */;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
output 	read_latency_shift_reg_0;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
output 	av_readdata_pre_6;
output 	av_readdata_pre_7;
input 	reset;
input 	write;
input 	write1;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter~0_combout ;
wire \wait_latency_counter~1_combout ;


dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(write1),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

cyclonev_lcell_comb \wait_latency_counter~0 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!write),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~0 .extended_lut = "off";
defparam \wait_latency_counter~0 .lut_mask = 64'h0404040404040404;
defparam \wait_latency_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(gnd),
	.datab(!wait_latency_counter_0),
	.datac(!write),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'h0C0C0C0C0C0C0C0C;
defparam \wait_latency_counter~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_slave_translator_14 (
	waitrequest_reset_override,
	out_valid_reg,
	mem_used_1,
	WideOr0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	read_latency_shift_reg_0,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	reset,
	m0_write,
	cp_ready,
	in_data_reg_69,
	av_readdata,
	clk)/* synthesis synthesis_greybox=0 */;
input 	waitrequest_reset_override;
input 	out_valid_reg;
input 	mem_used_1;
input 	WideOr0;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
output 	read_latency_shift_reg_0;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
output 	av_readdata_pre_6;
input 	reset;
input 	m0_write;
input 	cp_ready;
input 	in_data_reg_69;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~0_combout ;
wire \wait_latency_counter[0]~0_combout ;
wire \wait_latency_counter~1_combout ;
wire \wait_latency_counter~2_combout ;
wire \read_latency_shift_reg~1_combout ;


dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!mem_used_1),
	.datab(!WideOr0),
	.datac(!out_valid_reg),
	.datad(!in_data_reg_69),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'h0002000200020002;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter[0]~0 (
	.dataa(!waitrequest_reset_override),
	.datab(!wait_latency_counter_1),
	.datac(!wait_latency_counter_0),
	.datad(!m0_write),
	.datae(!\read_latency_shift_reg~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter[0]~0 .extended_lut = "off";
defparam \wait_latency_counter[0]~0 .lut_mask = 64'h0015511500155115;
defparam \wait_latency_counter[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!\wait_latency_counter[0]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'h0606060606060606;
defparam \wait_latency_counter~1 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~2 (
	.dataa(!wait_latency_counter_0),
	.datab(!\wait_latency_counter[0]~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~2 .extended_lut = "off";
defparam \wait_latency_counter~2 .lut_mask = 64'h2222222222222222;
defparam \wait_latency_counter~2 .shared_arith = "off";

cyclonev_lcell_comb \read_latency_shift_reg~1 (
	.dataa(!cp_ready),
	.datab(!\read_latency_shift_reg~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~1 .extended_lut = "off";
defparam \read_latency_shift_reg~1 .lut_mask = 64'h1111111111111111;
defparam \read_latency_shift_reg~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_slave_translator_15 (
	wait_latency_counter_1,
	wait_latency_counter_0,
	read_latency_shift_reg_0,
	av_readdata_pre_0,
	reset,
	write,
	write1,
	av_readdata,
	clk)/* synthesis synthesis_greybox=0 */;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
output 	read_latency_shift_reg_0;
output 	av_readdata_pre_0;
input 	reset;
input 	write;
input 	write1;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter~0_combout ;
wire \wait_latency_counter~1_combout ;


dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(write1),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

cyclonev_lcell_comb \wait_latency_counter~0 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!write),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~0 .extended_lut = "off";
defparam \wait_latency_counter~0 .lut_mask = 64'h0404040404040404;
defparam \wait_latency_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(gnd),
	.datab(!wait_latency_counter_0),
	.datac(!write),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'h0C0C0C0C0C0C0C0C;
defparam \wait_latency_counter~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_slave_translator_16 (
	waitrequest_reset_override,
	out_valid_reg,
	mem_used_1,
	WideOr0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	read_latency_shift_reg_0,
	av_readdata_pre_0,
	reset,
	m0_write,
	cp_ready,
	in_data_reg_69,
	av_readdata,
	clk)/* synthesis synthesis_greybox=0 */;
input 	waitrequest_reset_override;
input 	out_valid_reg;
input 	mem_used_1;
input 	WideOr0;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
output 	read_latency_shift_reg_0;
output 	av_readdata_pre_0;
input 	reset;
input 	m0_write;
input 	cp_ready;
input 	in_data_reg_69;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~0_combout ;
wire \wait_latency_counter[1]~0_combout ;
wire \wait_latency_counter~1_combout ;
wire \wait_latency_counter~2_combout ;
wire \read_latency_shift_reg~1_combout ;


dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!mem_used_1),
	.datab(!WideOr0),
	.datac(!out_valid_reg),
	.datad(!in_data_reg_69),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'h0002000200020002;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter[1]~0 (
	.dataa(!waitrequest_reset_override),
	.datab(!wait_latency_counter_1),
	.datac(!wait_latency_counter_0),
	.datad(!m0_write),
	.datae(!\read_latency_shift_reg~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter[1]~0 .extended_lut = "off";
defparam \wait_latency_counter[1]~0 .lut_mask = 64'h0015511500155115;
defparam \wait_latency_counter[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!\wait_latency_counter[1]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'h0606060606060606;
defparam \wait_latency_counter~1 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~2 (
	.dataa(!wait_latency_counter_0),
	.datab(!\wait_latency_counter[1]~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~2 .extended_lut = "off";
defparam \wait_latency_counter~2 .lut_mask = 64'h2222222222222222;
defparam \wait_latency_counter~2 .shared_arith = "off";

cyclonev_lcell_comb \read_latency_shift_reg~1 (
	.dataa(!cp_ready),
	.datab(!\read_latency_shift_reg~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~1 .extended_lut = "off";
defparam \read_latency_shift_reg~1 .lut_mask = 64'h1111111111111111;
defparam \read_latency_shift_reg~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_traffic_limiter (
	h2f_ARVALID_0,
	h2f_RREADY_0,
	has_pending_responses1,
	cmd_sink_data,
	last_channel_6,
	cmd_sink_channel,
	WideOr0,
	WideOr01,
	WideOr02,
	WideOr03,
	cmd_sink_ready,
	src_payload,
	src_payload_0,
	src_payload_01,
	src_payload_02,
	WideOr1,
	reset,
	last_channel_8,
	last_channel_11,
	last_channel_12,
	last_channel_1,
	last_channel_15,
	last_channel_16,
	last_channel_13,
	last_channel_14,
	last_channel_3,
	cmd_src_valid_5,
	last_channel_9,
	last_channel_10,
	last_channel_0,
	last_channel_4,
	last_channel_7,
	last_channel_2,
	clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARVALID_0;
input 	h2f_RREADY_0;
output 	has_pending_responses1;
input 	[128:0] cmd_sink_data;
output 	last_channel_6;
input 	[16:0] cmd_sink_channel;
input 	WideOr0;
input 	WideOr01;
input 	WideOr02;
input 	WideOr03;
output 	cmd_sink_ready;
input 	src_payload;
input 	src_payload_0;
input 	src_payload_01;
input 	src_payload_02;
input 	WideOr1;
input 	reset;
output 	last_channel_8;
output 	last_channel_11;
output 	last_channel_12;
output 	last_channel_1;
output 	last_channel_15;
output 	last_channel_16;
output 	last_channel_13;
output 	last_channel_14;
output 	last_channel_3;
output 	cmd_src_valid_5;
output 	last_channel_9;
output 	last_channel_10;
output 	last_channel_0;
output 	last_channel_4;
output 	last_channel_7;
output 	last_channel_2;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \last_dest_id[2]~q ;
wire \Equal0~0_combout ;
wire \last_dest_id[0]~q ;
wire \last_dest_id[1]~q ;
wire \last_dest_id[3]~q ;
wire \Equal0~1_combout ;
wire \save_dest_id~0_combout ;
wire \nonposted_cmd_accepted~combout ;
wire \pending_response_count[0]~1_combout ;
wire \response_sink_accepted~combout ;
wire \pending_response_count[1]~0_combout ;
wire \pending_response_count[0]~q ;
wire \Add0~0_combout ;
wire \pending_response_count[1]~q ;
wire \has_pending_responses~0_combout ;
wire \suppress_change_dest_id~combout ;
wire \last_channel[5]~q ;


dffeas has_pending_responses(
	.clk(clk),
	.d(\has_pending_responses~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(has_pending_responses1),
	.prn(vcc));
defparam has_pending_responses.is_wysiwyg = "true";
defparam has_pending_responses.power_up = "low";

dffeas \last_channel[6] (
	.clk(clk),
	.d(cmd_sink_channel[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(last_channel_6),
	.prn(vcc));
defparam \last_channel[6] .is_wysiwyg = "true";
defparam \last_channel[6] .power_up = "low";

cyclonev_lcell_comb \cmd_sink_ready~0 (
	.dataa(!\suppress_change_dest_id~combout ),
	.datab(!WideOr0),
	.datac(!WideOr01),
	.datad(!WideOr02),
	.datae(!WideOr03),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cmd_sink_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \cmd_sink_ready~0 .extended_lut = "off";
defparam \cmd_sink_ready~0 .lut_mask = 64'hAAAAAAA8AAAAAAA8;
defparam \cmd_sink_ready~0 .shared_arith = "off";

dffeas \last_channel[8] (
	.clk(clk),
	.d(cmd_sink_channel[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(last_channel_8),
	.prn(vcc));
defparam \last_channel[8] .is_wysiwyg = "true";
defparam \last_channel[8] .power_up = "low";

dffeas \last_channel[11] (
	.clk(clk),
	.d(cmd_sink_channel[11]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(last_channel_11),
	.prn(vcc));
defparam \last_channel[11] .is_wysiwyg = "true";
defparam \last_channel[11] .power_up = "low";

dffeas \last_channel[12] (
	.clk(clk),
	.d(cmd_sink_channel[12]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(last_channel_12),
	.prn(vcc));
defparam \last_channel[12] .is_wysiwyg = "true";
defparam \last_channel[12] .power_up = "low";

dffeas \last_channel[1] (
	.clk(clk),
	.d(cmd_sink_channel[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(last_channel_1),
	.prn(vcc));
defparam \last_channel[1] .is_wysiwyg = "true";
defparam \last_channel[1] .power_up = "low";

dffeas \last_channel[15] (
	.clk(clk),
	.d(cmd_sink_channel[15]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(last_channel_15),
	.prn(vcc));
defparam \last_channel[15] .is_wysiwyg = "true";
defparam \last_channel[15] .power_up = "low";

dffeas \last_channel[16] (
	.clk(clk),
	.d(cmd_sink_channel[16]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(last_channel_16),
	.prn(vcc));
defparam \last_channel[16] .is_wysiwyg = "true";
defparam \last_channel[16] .power_up = "low";

dffeas \last_channel[13] (
	.clk(clk),
	.d(cmd_sink_channel[13]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(last_channel_13),
	.prn(vcc));
defparam \last_channel[13] .is_wysiwyg = "true";
defparam \last_channel[13] .power_up = "low";

dffeas \last_channel[14] (
	.clk(clk),
	.d(cmd_sink_channel[14]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(last_channel_14),
	.prn(vcc));
defparam \last_channel[14] .is_wysiwyg = "true";
defparam \last_channel[14] .power_up = "low";

dffeas \last_channel[3] (
	.clk(clk),
	.d(cmd_sink_channel[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(last_channel_3),
	.prn(vcc));
defparam \last_channel[3] .is_wysiwyg = "true";
defparam \last_channel[3] .power_up = "low";

cyclonev_lcell_comb \cmd_src_valid[5]~0 (
	.dataa(!has_pending_responses1),
	.datab(!\last_channel[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cmd_src_valid_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \cmd_src_valid[5]~0 .extended_lut = "off";
defparam \cmd_src_valid[5]~0 .lut_mask = 64'h4444444444444444;
defparam \cmd_src_valid[5]~0 .shared_arith = "off";

dffeas \last_channel[9] (
	.clk(clk),
	.d(cmd_sink_channel[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(last_channel_9),
	.prn(vcc));
defparam \last_channel[9] .is_wysiwyg = "true";
defparam \last_channel[9] .power_up = "low";

dffeas \last_channel[10] (
	.clk(clk),
	.d(cmd_sink_channel[10]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(last_channel_10),
	.prn(vcc));
defparam \last_channel[10] .is_wysiwyg = "true";
defparam \last_channel[10] .power_up = "low";

dffeas \last_channel[0] (
	.clk(clk),
	.d(cmd_sink_channel[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(last_channel_0),
	.prn(vcc));
defparam \last_channel[0] .is_wysiwyg = "true";
defparam \last_channel[0] .power_up = "low";

dffeas \last_channel[4] (
	.clk(clk),
	.d(cmd_sink_channel[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(last_channel_4),
	.prn(vcc));
defparam \last_channel[4] .is_wysiwyg = "true";
defparam \last_channel[4] .power_up = "low";

dffeas \last_channel[7] (
	.clk(clk),
	.d(cmd_sink_channel[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(last_channel_7),
	.prn(vcc));
defparam \last_channel[7] .is_wysiwyg = "true";
defparam \last_channel[7] .power_up = "low";

dffeas \last_channel[2] (
	.clk(clk),
	.d(cmd_sink_channel[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(last_channel_2),
	.prn(vcc));
defparam \last_channel[2] .is_wysiwyg = "true";
defparam \last_channel[2] .power_up = "low";

dffeas \last_dest_id[2] (
	.clk(clk),
	.d(cmd_sink_data[102]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(\last_dest_id[2]~q ),
	.prn(vcc));
defparam \last_dest_id[2] .is_wysiwyg = "true";
defparam \last_dest_id[2] .power_up = "low";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!\last_dest_id[2]~q ),
	.datab(!cmd_sink_data[102]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'h6666666666666666;
defparam \Equal0~0 .shared_arith = "off";

dffeas \last_dest_id[0] (
	.clk(clk),
	.d(cmd_sink_data[100]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(\last_dest_id[0]~q ),
	.prn(vcc));
defparam \last_dest_id[0] .is_wysiwyg = "true";
defparam \last_dest_id[0] .power_up = "low";

dffeas \last_dest_id[1] (
	.clk(clk),
	.d(cmd_sink_data[101]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(\last_dest_id[1]~q ),
	.prn(vcc));
defparam \last_dest_id[1] .is_wysiwyg = "true";
defparam \last_dest_id[1] .power_up = "low";

dffeas \last_dest_id[3] (
	.clk(clk),
	.d(cmd_sink_data[103]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(\last_dest_id[3]~q ),
	.prn(vcc));
defparam \last_dest_id[3] .is_wysiwyg = "true";
defparam \last_dest_id[3] .power_up = "low";

cyclonev_lcell_comb \Equal0~1 (
	.dataa(!\last_dest_id[0]~q ),
	.datab(!cmd_sink_data[100]),
	.datac(!\last_dest_id[1]~q ),
	.datad(!cmd_sink_data[101]),
	.datae(!\last_dest_id[3]~q ),
	.dataf(!cmd_sink_data[103]),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~1 .extended_lut = "off";
defparam \Equal0~1 .lut_mask = 64'h9009000000009009;
defparam \Equal0~1 .shared_arith = "off";

cyclonev_lcell_comb \save_dest_id~0 (
	.dataa(!h2f_ARVALID_0),
	.datab(!has_pending_responses1),
	.datac(!\Equal0~0_combout ),
	.datad(!last_channel_6),
	.datae(!cmd_sink_channel[6]),
	.dataf(!\Equal0~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\save_dest_id~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \save_dest_id~0 .extended_lut = "off";
defparam \save_dest_id~0 .lut_mask = 64'h4444444454444454;
defparam \save_dest_id~0 .shared_arith = "off";

cyclonev_lcell_comb nonposted_cmd_accepted(
	.dataa(!WideOr0),
	.datab(!WideOr01),
	.datac(!WideOr02),
	.datad(!WideOr03),
	.datae(!\save_dest_id~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nonposted_cmd_accepted~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam nonposted_cmd_accepted.extended_lut = "off";
defparam nonposted_cmd_accepted.lut_mask = 64'h0000FFFE0000FFFE;
defparam nonposted_cmd_accepted.shared_arith = "off";

cyclonev_lcell_comb \pending_response_count[0]~1 (
	.dataa(!\pending_response_count[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pending_response_count[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pending_response_count[0]~1 .extended_lut = "off";
defparam \pending_response_count[0]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \pending_response_count[0]~1 .shared_arith = "off";

cyclonev_lcell_comb response_sink_accepted(
	.dataa(!h2f_RREADY_0),
	.datab(!src_payload),
	.datac(!src_payload_0),
	.datad(!src_payload_01),
	.datae(!src_payload_02),
	.dataf(!WideOr1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\response_sink_accepted~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam response_sink_accepted.extended_lut = "off";
defparam response_sink_accepted.lut_mask = 64'h0000000055555551;
defparam response_sink_accepted.shared_arith = "off";

cyclonev_lcell_comb \pending_response_count[1]~0 (
	.dataa(!WideOr0),
	.datab(!WideOr01),
	.datac(!WideOr02),
	.datad(!WideOr03),
	.datae(!\save_dest_id~0_combout ),
	.dataf(!\response_sink_accepted~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pending_response_count[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pending_response_count[1]~0 .extended_lut = "off";
defparam \pending_response_count[1]~0 .lut_mask = 64'h0000FFFEFFFF0001;
defparam \pending_response_count[1]~0 .shared_arith = "off";

dffeas \pending_response_count[0] (
	.clk(clk),
	.d(\pending_response_count[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pending_response_count[1]~0_combout ),
	.q(\pending_response_count[0]~q ),
	.prn(vcc));
defparam \pending_response_count[0] .is_wysiwyg = "true";
defparam \pending_response_count[0] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!\pending_response_count[1]~q ),
	.datab(!\pending_response_count[0]~q ),
	.datac(!\response_sink_accepted~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h6969696969696969;
defparam \Add0~0 .shared_arith = "off";

dffeas \pending_response_count[1] (
	.clk(clk),
	.d(\Add0~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pending_response_count[1]~0_combout ),
	.q(\pending_response_count[1]~q ),
	.prn(vcc));
defparam \pending_response_count[1] .is_wysiwyg = "true";
defparam \pending_response_count[1] .power_up = "low";

cyclonev_lcell_comb \has_pending_responses~0 (
	.dataa(!has_pending_responses1),
	.datab(!\nonposted_cmd_accepted~combout ),
	.datac(!\pending_response_count[1]~q ),
	.datad(!\pending_response_count[0]~q ),
	.datae(!\response_sink_accepted~combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\has_pending_responses~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \has_pending_responses~0 .extended_lut = "off";
defparam \has_pending_responses~0 .lut_mask = 64'h7555551575555515;
defparam \has_pending_responses~0 .shared_arith = "off";

cyclonev_lcell_comb suppress_change_dest_id(
	.dataa(!has_pending_responses1),
	.datab(!\Equal0~0_combout ),
	.datac(!last_channel_6),
	.datad(!cmd_sink_channel[6]),
	.datae(!\Equal0~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\suppress_change_dest_id~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam suppress_change_dest_id.extended_lut = "off";
defparam suppress_change_dest_id.lut_mask = 64'h5555155155551551;
defparam suppress_change_dest_id.shared_arith = "off";

dffeas \last_channel[5] (
	.clk(clk),
	.d(cmd_sink_channel[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(\last_channel[5]~q ),
	.prn(vcc));
defparam \last_channel[5] .is_wysiwyg = "true";
defparam \last_channel[5] .power_up = "low";

endmodule

module spw_babasu_altera_merlin_traffic_limiter_1 (
	h2f_BREADY_0,
	h2f_WLAST_0,
	write_addr_data_both_valid,
	has_pending_responses1,
	out_data_4,
	cmd_sink_data,
	Equal5,
	Equal14,
	last_channel_6,
	WideOr0,
	WideOr01,
	WideOr02,
	WideOr03,
	WideOr04,
	WideOr05,
	nonposted_cmd_accepted,
	WideOr1,
	nonposted_cmd_accepted1,
	reset,
	last_channel_1,
	last_channel_15,
	last_channel_16,
	last_channel_13,
	last_channel_14,
	last_channel_5,
	last_channel_9,
	last_channel_0,
	last_channel_2,
	src_payload,
	src_payload1,
	src_payload_0,
	src_payload_01,
	cmd_sink_channel,
	clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_BREADY_0;
input 	h2f_WLAST_0;
input 	write_addr_data_both_valid;
output 	has_pending_responses1;
input 	out_data_4;
input 	[128:0] cmd_sink_data;
input 	Equal5;
input 	Equal14;
output 	last_channel_6;
input 	WideOr0;
input 	WideOr01;
input 	WideOr02;
input 	WideOr03;
input 	WideOr04;
input 	WideOr05;
output 	nonposted_cmd_accepted;
input 	WideOr1;
output 	nonposted_cmd_accepted1;
input 	reset;
output 	last_channel_1;
output 	last_channel_15;
output 	last_channel_16;
output 	last_channel_13;
output 	last_channel_14;
output 	last_channel_5;
output 	last_channel_9;
output 	last_channel_0;
output 	last_channel_2;
input 	src_payload;
input 	src_payload1;
input 	src_payload_0;
input 	src_payload_01;
input 	[16:0] cmd_sink_channel;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \last_dest_id[2]~q ;
wire \Equal0~0_combout ;
wire \last_dest_id[0]~q ;
wire \last_dest_id[1]~q ;
wire \last_dest_id[3]~q ;
wire \Equal0~1_combout ;
wire \save_dest_id~0_combout ;
wire \pending_response_count[0]~1_combout ;
wire \response_sink_accepted~combout ;
wire \pending_response_count[1]~0_combout ;
wire \pending_response_count[0]~q ;
wire \Add0~0_combout ;
wire \pending_response_count[1]~q ;
wire \has_pending_responses~0_combout ;
wire \has_pending_responses~1_combout ;
wire \has_pending_responses~2_combout ;


dffeas has_pending_responses(
	.clk(clk),
	.d(\has_pending_responses~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(has_pending_responses1),
	.prn(vcc));
defparam has_pending_responses.is_wysiwyg = "true";
defparam has_pending_responses.power_up = "low";

dffeas \last_channel[6] (
	.clk(clk),
	.d(cmd_sink_channel[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(last_channel_6),
	.prn(vcc));
defparam \last_channel[6] .is_wysiwyg = "true";
defparam \last_channel[6] .power_up = "low";

cyclonev_lcell_comb \nonposted_cmd_accepted~0 (
	.dataa(!h2f_WLAST_0),
	.datab(!\save_dest_id~0_combout ),
	.datac(!WideOr0),
	.datad(!WideOr05),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nonposted_cmd_accepted),
	.sumout(),
	.cout(),
	.shareout());
defparam \nonposted_cmd_accepted~0 .extended_lut = "off";
defparam \nonposted_cmd_accepted~0 .lut_mask = 64'h1110111011101110;
defparam \nonposted_cmd_accepted~0 .shared_arith = "off";

cyclonev_lcell_comb \nonposted_cmd_accepted~1 (
	.dataa(!\save_dest_id~0_combout ),
	.datab(!WideOr0),
	.datac(!WideOr01),
	.datad(!WideOr02),
	.datae(!WideOr03),
	.dataf(!WideOr04),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nonposted_cmd_accepted1),
	.sumout(),
	.cout(),
	.shareout());
defparam \nonposted_cmd_accepted~1 .extended_lut = "off";
defparam \nonposted_cmd_accepted~1 .lut_mask = 64'h5555555555555554;
defparam \nonposted_cmd_accepted~1 .shared_arith = "off";

dffeas \last_channel[1] (
	.clk(clk),
	.d(cmd_sink_channel[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(last_channel_1),
	.prn(vcc));
defparam \last_channel[1] .is_wysiwyg = "true";
defparam \last_channel[1] .power_up = "low";

dffeas \last_channel[15] (
	.clk(clk),
	.d(cmd_sink_channel[15]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(last_channel_15),
	.prn(vcc));
defparam \last_channel[15] .is_wysiwyg = "true";
defparam \last_channel[15] .power_up = "low";

dffeas \last_channel[16] (
	.clk(clk),
	.d(cmd_sink_channel[16]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(last_channel_16),
	.prn(vcc));
defparam \last_channel[16] .is_wysiwyg = "true";
defparam \last_channel[16] .power_up = "low";

dffeas \last_channel[13] (
	.clk(clk),
	.d(cmd_sink_channel[13]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(last_channel_13),
	.prn(vcc));
defparam \last_channel[13] .is_wysiwyg = "true";
defparam \last_channel[13] .power_up = "low";

dffeas \last_channel[14] (
	.clk(clk),
	.d(cmd_sink_channel[14]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(last_channel_14),
	.prn(vcc));
defparam \last_channel[14] .is_wysiwyg = "true";
defparam \last_channel[14] .power_up = "low";

dffeas \last_channel[5] (
	.clk(clk),
	.d(cmd_sink_channel[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(last_channel_5),
	.prn(vcc));
defparam \last_channel[5] .is_wysiwyg = "true";
defparam \last_channel[5] .power_up = "low";

dffeas \last_channel[9] (
	.clk(clk),
	.d(cmd_sink_channel[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(last_channel_9),
	.prn(vcc));
defparam \last_channel[9] .is_wysiwyg = "true";
defparam \last_channel[9] .power_up = "low";

dffeas \last_channel[0] (
	.clk(clk),
	.d(cmd_sink_channel[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(last_channel_0),
	.prn(vcc));
defparam \last_channel[0] .is_wysiwyg = "true";
defparam \last_channel[0] .power_up = "low";

dffeas \last_channel[2] (
	.clk(clk),
	.d(cmd_sink_channel[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(last_channel_2),
	.prn(vcc));
defparam \last_channel[2] .is_wysiwyg = "true";
defparam \last_channel[2] .power_up = "low";

dffeas \last_dest_id[2] (
	.clk(clk),
	.d(cmd_sink_data[102]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(\last_dest_id[2]~q ),
	.prn(vcc));
defparam \last_dest_id[2] .is_wysiwyg = "true";
defparam \last_dest_id[2] .power_up = "low";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!out_data_4),
	.datab(!Equal5),
	.datac(!Equal14),
	.datad(!last_channel_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'hFD02FD02FD02FD02;
defparam \Equal0~0 .shared_arith = "off";

dffeas \last_dest_id[0] (
	.clk(clk),
	.d(cmd_sink_data[100]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(\last_dest_id[0]~q ),
	.prn(vcc));
defparam \last_dest_id[0] .is_wysiwyg = "true";
defparam \last_dest_id[0] .power_up = "low";

dffeas \last_dest_id[1] (
	.clk(clk),
	.d(cmd_sink_data[101]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(\last_dest_id[1]~q ),
	.prn(vcc));
defparam \last_dest_id[1] .is_wysiwyg = "true";
defparam \last_dest_id[1] .power_up = "low";

dffeas \last_dest_id[3] (
	.clk(clk),
	.d(cmd_sink_data[103]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(\last_dest_id[3]~q ),
	.prn(vcc));
defparam \last_dest_id[3] .is_wysiwyg = "true";
defparam \last_dest_id[3] .power_up = "low";

cyclonev_lcell_comb \Equal0~1 (
	.dataa(!\last_dest_id[0]~q ),
	.datab(!cmd_sink_data[100]),
	.datac(!\last_dest_id[1]~q ),
	.datad(!cmd_sink_data[101]),
	.datae(!\last_dest_id[3]~q ),
	.dataf(!cmd_sink_data[103]),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~1 .extended_lut = "off";
defparam \Equal0~1 .lut_mask = 64'h9009000000009009;
defparam \Equal0~1 .shared_arith = "off";

cyclonev_lcell_comb \save_dest_id~0 (
	.dataa(!write_addr_data_both_valid),
	.datab(!has_pending_responses1),
	.datac(!\last_dest_id[2]~q ),
	.datad(!cmd_sink_data[102]),
	.datae(!\Equal0~0_combout ),
	.dataf(!\Equal0~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\save_dest_id~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \save_dest_id~0 .extended_lut = "off";
defparam \save_dest_id~0 .lut_mask = 64'h4444444444445445;
defparam \save_dest_id~0 .shared_arith = "off";

cyclonev_lcell_comb \pending_response_count[0]~1 (
	.dataa(!\pending_response_count[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pending_response_count[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pending_response_count[0]~1 .extended_lut = "off";
defparam \pending_response_count[0]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \pending_response_count[0]~1 .shared_arith = "off";

cyclonev_lcell_comb response_sink_accepted(
	.dataa(!h2f_BREADY_0),
	.datab(!src_payload),
	.datac(!src_payload1),
	.datad(!src_payload_0),
	.datae(!src_payload_01),
	.dataf(!WideOr1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\response_sink_accepted~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam response_sink_accepted.extended_lut = "off";
defparam response_sink_accepted.lut_mask = 64'h0000000055155555;
defparam response_sink_accepted.shared_arith = "off";

cyclonev_lcell_comb \pending_response_count[1]~0 (
	.dataa(!h2f_WLAST_0),
	.datab(!\save_dest_id~0_combout ),
	.datac(!WideOr0),
	.datad(!WideOr05),
	.datae(!\response_sink_accepted~combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pending_response_count[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pending_response_count[1]~0 .extended_lut = "off";
defparam \pending_response_count[1]~0 .lut_mask = 64'h1110EEEF1110EEEF;
defparam \pending_response_count[1]~0 .shared_arith = "off";

dffeas \pending_response_count[0] (
	.clk(clk),
	.d(\pending_response_count[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pending_response_count[1]~0_combout ),
	.q(\pending_response_count[0]~q ),
	.prn(vcc));
defparam \pending_response_count[0] .is_wysiwyg = "true";
defparam \pending_response_count[0] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!\pending_response_count[1]~q ),
	.datab(!\pending_response_count[0]~q ),
	.datac(!\response_sink_accepted~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h6969696969696969;
defparam \Add0~0 .shared_arith = "off";

dffeas \pending_response_count[1] (
	.clk(clk),
	.d(\Add0~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pending_response_count[1]~0_combout ),
	.q(\pending_response_count[1]~q ),
	.prn(vcc));
defparam \pending_response_count[1] .is_wysiwyg = "true";
defparam \pending_response_count[1] .power_up = "low";

cyclonev_lcell_comb \has_pending_responses~0 (
	.dataa(!has_pending_responses1),
	.datab(!\pending_response_count[1]~q ),
	.datac(!\pending_response_count[0]~q ),
	.datad(!\response_sink_accepted~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\has_pending_responses~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \has_pending_responses~0 .extended_lut = "off";
defparam \has_pending_responses~0 .lut_mask = 64'h2AAA2AAA2AAA2AAA;
defparam \has_pending_responses~0 .shared_arith = "off";

cyclonev_lcell_comb \has_pending_responses~1 (
	.dataa(!has_pending_responses1),
	.datab(!\pending_response_count[1]~q ),
	.datac(!\pending_response_count[0]~q ),
	.datad(!\response_sink_accepted~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\has_pending_responses~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \has_pending_responses~1 .extended_lut = "off";
defparam \has_pending_responses~1 .lut_mask = 64'h5551555155515551;
defparam \has_pending_responses~1 .shared_arith = "off";

cyclonev_lcell_comb \has_pending_responses~2 (
	.dataa(!h2f_WLAST_0),
	.datab(!\save_dest_id~0_combout ),
	.datac(!WideOr0),
	.datad(!WideOr05),
	.datae(!\has_pending_responses~0_combout ),
	.dataf(!\has_pending_responses~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\has_pending_responses~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \has_pending_responses~2 .extended_lut = "off";
defparam \has_pending_responses~2 .lut_mask = 64'h11100000FFFFFFFF;
defparam \has_pending_responses~2 .shared_arith = "off";

endmodule

module spw_babasu_spw_babasu_mm_interconnect_0_cmd_demux (
	h2f_AWVALID_0,
	h2f_WVALID_0,
	nxt_in_ready,
	nxt_in_ready1,
	nxt_in_ready2,
	nxt_in_ready3,
	nxt_in_ready4,
	nxt_in_ready5,
	nxt_in_ready6,
	nxt_in_ready7,
	nxt_in_ready8,
	nxt_in_ready9,
	nxt_in_ready10,
	nxt_in_ready11,
	nxt_in_ready12,
	nxt_in_ready13,
	nxt_in_ready14,
	nxt_in_ready15,
	nxt_in_ready16,
	nxt_in_ready17,
	nxt_in_ready18,
	nxt_in_ready19,
	write_addr_data_both_valid,
	has_pending_responses,
	out_data_8,
	out_data_5,
	out_data_4,
	out_data_7,
	out_data_6,
	Equal5,
	Equal14,
	last_channel_6,
	Equal16,
	Equal13,
	Equal15,
	saved_grant_0,
	Equal161,
	saved_grant_01,
	WideOr0,
	saved_grant_02,
	saved_grant_03,
	WideOr01,
	saved_grant_04,
	Equal9,
	saved_grant_05,
	WideOr02,
	saved_grant_06,
	saved_grant_07,
	WideOr03,
	saved_grant_08,
	saved_grant_09,
	WideOr04,
	WideOr05,
	last_channel_1,
	src1_valid,
	src1_valid1,
	src1_valid2,
	last_channel_15,
	src15_valid,
	src15_valid1,
	src15_valid2,
	last_channel_16,
	src16_valid,
	src16_valid1,
	src16_valid2,
	last_channel_13,
	src13_valid,
	src13_valid1,
	src13_valid2,
	last_channel_14,
	src14_valid,
	src14_valid1,
	src14_valid2,
	last_channel_5,
	src5_valid,
	src5_valid1,
	src5_valid2,
	last_channel_9,
	src9_valid,
	src9_valid1,
	src9_valid2,
	last_channel_0,
	src0_valid,
	last_channel_2,
	src2_valid,
	src2_valid1,
	src2_valid2,
	src6_valid,
	src6_valid1,
	src6_valid2)/* synthesis synthesis_greybox=0 */;
input 	h2f_AWVALID_0;
input 	h2f_WVALID_0;
input 	nxt_in_ready;
input 	nxt_in_ready1;
input 	nxt_in_ready2;
input 	nxt_in_ready3;
input 	nxt_in_ready4;
input 	nxt_in_ready5;
input 	nxt_in_ready6;
input 	nxt_in_ready7;
input 	nxt_in_ready8;
input 	nxt_in_ready9;
input 	nxt_in_ready10;
input 	nxt_in_ready11;
input 	nxt_in_ready12;
input 	nxt_in_ready13;
input 	nxt_in_ready14;
input 	nxt_in_ready15;
input 	nxt_in_ready16;
input 	nxt_in_ready17;
input 	nxt_in_ready18;
input 	nxt_in_ready19;
input 	write_addr_data_both_valid;
input 	has_pending_responses;
input 	out_data_8;
input 	out_data_5;
input 	out_data_4;
input 	out_data_7;
input 	out_data_6;
input 	Equal5;
input 	Equal14;
input 	last_channel_6;
input 	Equal16;
input 	Equal13;
input 	Equal15;
input 	saved_grant_0;
input 	Equal161;
input 	saved_grant_01;
output 	WideOr0;
input 	saved_grant_02;
input 	saved_grant_03;
output 	WideOr01;
input 	saved_grant_04;
input 	Equal9;
input 	saved_grant_05;
output 	WideOr02;
input 	saved_grant_06;
input 	saved_grant_07;
output 	WideOr03;
input 	saved_grant_08;
input 	saved_grant_09;
output 	WideOr04;
output 	WideOr05;
input 	last_channel_1;
output 	src1_valid;
output 	src1_valid1;
output 	src1_valid2;
input 	last_channel_15;
output 	src15_valid;
output 	src15_valid1;
output 	src15_valid2;
input 	last_channel_16;
output 	src16_valid;
output 	src16_valid1;
output 	src16_valid2;
input 	last_channel_13;
output 	src13_valid;
output 	src13_valid1;
output 	src13_valid2;
input 	last_channel_14;
output 	src14_valid;
output 	src14_valid1;
output 	src14_valid2;
input 	last_channel_5;
output 	src5_valid;
output 	src5_valid1;
output 	src5_valid2;
input 	last_channel_9;
output 	src9_valid;
output 	src9_valid1;
output 	src9_valid2;
input 	last_channel_0;
output 	src0_valid;
input 	last_channel_2;
output 	src2_valid;
output 	src2_valid1;
output 	src2_valid2;
output 	src6_valid;
output 	src6_valid1;
output 	src6_valid2;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \sink_ready~0_combout ;
wire \sink_ready~1_combout ;
wire \sink_ready~2_combout ;
wire \sink_ready~3_combout ;
wire \sink_ready~4_combout ;
wire \sink_ready~5_combout ;
wire \sink_ready~6_combout ;
wire \sink_ready~7_combout ;
wire \sink_ready~8_combout ;
wire \sink_ready~9_combout ;
wire \src0_valid~0_combout ;


cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!nxt_in_ready11),
	.datab(!nxt_in_ready8),
	.datac(!nxt_in_ready12),
	.datad(!nxt_in_ready7),
	.datae(!\sink_ready~0_combout ),
	.dataf(!\sink_ready~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'hFFFF8888F0008000;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~1 (
	.dataa(!nxt_in_ready13),
	.datab(!nxt_in_ready6),
	.datac(!nxt_in_ready14),
	.datad(!nxt_in_ready5),
	.datae(!\sink_ready~2_combout ),
	.dataf(!\sink_ready~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr01),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~1 .extended_lut = "off";
defparam \WideOr0~1 .lut_mask = 64'hFFFF8888F0008000;
defparam \WideOr0~1 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~2 (
	.dataa(!nxt_in_ready16),
	.datab(!nxt_in_ready3),
	.datac(!nxt_in_ready19),
	.datad(!nxt_in_ready),
	.datae(!\sink_ready~4_combout ),
	.dataf(!\sink_ready~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr02),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~2 .extended_lut = "off";
defparam \WideOr0~2 .lut_mask = 64'hFFFFF00088888000;
defparam \WideOr0~2 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~3 (
	.dataa(!nxt_in_ready10),
	.datab(!nxt_in_ready9),
	.datac(!nxt_in_ready17),
	.datad(!nxt_in_ready2),
	.datae(!\sink_ready~6_combout ),
	.dataf(!\sink_ready~7_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr03),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~3 .extended_lut = "off";
defparam \WideOr0~3 .lut_mask = 64'hFFFFF00088888000;
defparam \WideOr0~3 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~4 (
	.dataa(!nxt_in_ready15),
	.datab(!nxt_in_ready4),
	.datac(!nxt_in_ready18),
	.datad(!nxt_in_ready1),
	.datae(!\sink_ready~8_combout ),
	.dataf(!\sink_ready~9_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr04),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~4 .extended_lut = "off";
defparam \WideOr0~4 .lut_mask = 64'hFFFFF00088888000;
defparam \WideOr0~4 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~5 (
	.dataa(!WideOr01),
	.datab(!WideOr02),
	.datac(!WideOr03),
	.datad(!WideOr04),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr05),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~5 .extended_lut = "off";
defparam \WideOr0~5 .lut_mask = 64'h0001000100010001;
defparam \WideOr0~5 .shared_arith = "off";

cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!has_pending_responses),
	.datab(!last_channel_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'h4444444444444444;
defparam \src1_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src1_valid~1 (
	.dataa(!write_addr_data_both_valid),
	.datab(!src1_valid),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~1 .extended_lut = "off";
defparam \src1_valid~1 .lut_mask = 64'h4444444444444444;
defparam \src1_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \src1_valid~2 (
	.dataa(!out_data_5),
	.datab(!Equal16),
	.datac(!Equal15),
	.datad(!write_addr_data_both_valid),
	.datae(!src1_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~2 .extended_lut = "off";
defparam \src1_valid~2 .lut_mask = 64'h0002000000020000;
defparam \src1_valid~2 .shared_arith = "off";

cyclonev_lcell_comb \src15_valid~0 (
	.dataa(!has_pending_responses),
	.datab(!last_channel_15),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src15_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src15_valid~0 .extended_lut = "off";
defparam \src15_valid~0 .lut_mask = 64'h4444444444444444;
defparam \src15_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src15_valid~1 (
	.dataa(!write_addr_data_both_valid),
	.datab(!src15_valid),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src15_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src15_valid~1 .extended_lut = "off";
defparam \src15_valid~1 .lut_mask = 64'h4444444444444444;
defparam \src15_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \src15_valid~2 (
	.dataa(!out_data_5),
	.datab(!Equal15),
	.datac(!Equal13),
	.datad(!write_addr_data_both_valid),
	.datae(!src15_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src15_valid2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src15_valid~2 .extended_lut = "off";
defparam \src15_valid~2 .lut_mask = 64'h0001000000010000;
defparam \src15_valid~2 .shared_arith = "off";

cyclonev_lcell_comb \src16_valid~0 (
	.dataa(!has_pending_responses),
	.datab(!last_channel_16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src16_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src16_valid~0 .extended_lut = "off";
defparam \src16_valid~0 .lut_mask = 64'h4444444444444444;
defparam \src16_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src16_valid~1 (
	.dataa(!out_data_4),
	.datab(!Equal16),
	.datac(!Equal161),
	.datad(!write_addr_data_both_valid),
	.datae(!src16_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src16_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src16_valid~1 .extended_lut = "off";
defparam \src16_valid~1 .lut_mask = 64'h0002000000020000;
defparam \src16_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \src16_valid~2 (
	.dataa(!write_addr_data_both_valid),
	.datab(!src16_valid),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src16_valid2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src16_valid~2 .extended_lut = "off";
defparam \src16_valid~2 .lut_mask = 64'h4444444444444444;
defparam \src16_valid~2 .shared_arith = "off";

cyclonev_lcell_comb \src13_valid~0 (
	.dataa(!has_pending_responses),
	.datab(!last_channel_13),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src13_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src13_valid~0 .extended_lut = "off";
defparam \src13_valid~0 .lut_mask = 64'h4444444444444444;
defparam \src13_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src13_valid~1 (
	.dataa(!write_addr_data_both_valid),
	.datab(!src13_valid),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src13_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src13_valid~1 .extended_lut = "off";
defparam \src13_valid~1 .lut_mask = 64'h4444444444444444;
defparam \src13_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \src13_valid~2 (
	.dataa(!out_data_5),
	.datab(!Equal15),
	.datac(!Equal13),
	.datad(!write_addr_data_both_valid),
	.datae(!src13_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src13_valid2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src13_valid~2 .extended_lut = "off";
defparam \src13_valid~2 .lut_mask = 64'h0002000000020000;
defparam \src13_valid~2 .shared_arith = "off";

cyclonev_lcell_comb \src14_valid~0 (
	.dataa(!has_pending_responses),
	.datab(!last_channel_14),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src14_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src14_valid~0 .extended_lut = "off";
defparam \src14_valid~0 .lut_mask = 64'h4444444444444444;
defparam \src14_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src14_valid~1 (
	.dataa(!write_addr_data_both_valid),
	.datab(!src14_valid),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src14_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src14_valid~1 .extended_lut = "off";
defparam \src14_valid~1 .lut_mask = 64'h4444444444444444;
defparam \src14_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \src14_valid~2 (
	.dataa(!out_data_4),
	.datab(!Equal14),
	.datac(!Equal13),
	.datad(!write_addr_data_both_valid),
	.datae(!src14_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src14_valid2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src14_valid~2 .extended_lut = "off";
defparam \src14_valid~2 .lut_mask = 64'h0002000000020000;
defparam \src14_valid~2 .shared_arith = "off";

cyclonev_lcell_comb \src5_valid~0 (
	.dataa(!has_pending_responses),
	.datab(!last_channel_5),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src5_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src5_valid~0 .extended_lut = "off";
defparam \src5_valid~0 .lut_mask = 64'h4444444444444444;
defparam \src5_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src5_valid~1 (
	.dataa(!write_addr_data_both_valid),
	.datab(!src5_valid),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src5_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src5_valid~1 .extended_lut = "off";
defparam \src5_valid~1 .lut_mask = 64'h4444444444444444;
defparam \src5_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \src5_valid~2 (
	.dataa(!out_data_5),
	.datab(!Equal15),
	.datac(!Equal5),
	.datad(!write_addr_data_both_valid),
	.datae(!src5_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src5_valid2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src5_valid~2 .extended_lut = "off";
defparam \src5_valid~2 .lut_mask = 64'h0002000000020000;
defparam \src5_valid~2 .shared_arith = "off";

cyclonev_lcell_comb \src9_valid~0 (
	.dataa(!has_pending_responses),
	.datab(!last_channel_9),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src9_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src9_valid~0 .extended_lut = "off";
defparam \src9_valid~0 .lut_mask = 64'h4444444444444444;
defparam \src9_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src9_valid~1 (
	.dataa(!write_addr_data_both_valid),
	.datab(!src9_valid),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src9_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src9_valid~1 .extended_lut = "off";
defparam \src9_valid~1 .lut_mask = 64'h4444444444444444;
defparam \src9_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \src9_valid~2 (
	.dataa(!out_data_5),
	.datab(!Equal15),
	.datac(!Equal9),
	.datad(!write_addr_data_both_valid),
	.datae(!src9_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src9_valid2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src9_valid~2 .extended_lut = "off";
defparam \src9_valid~2 .lut_mask = 64'h0002000000020000;
defparam \src9_valid~2 .shared_arith = "off";

cyclonev_lcell_comb \src0_valid~1 (
	.dataa(!out_data_8),
	.datab(!out_data_5),
	.datac(!out_data_4),
	.datad(!out_data_7),
	.datae(!out_data_6),
	.dataf(!\src0_valid~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src0_valid~1 .extended_lut = "off";
defparam \src0_valid~1 .lut_mask = 64'h0000000097F7D7D5;
defparam \src0_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \src2_valid~0 (
	.dataa(!has_pending_responses),
	.datab(!last_channel_2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src2_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src2_valid~0 .extended_lut = "off";
defparam \src2_valid~0 .lut_mask = 64'h4444444444444444;
defparam \src2_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src2_valid~1 (
	.dataa(!write_addr_data_both_valid),
	.datab(!src2_valid),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src2_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src2_valid~1 .extended_lut = "off";
defparam \src2_valid~1 .lut_mask = 64'h4444444444444444;
defparam \src2_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \src2_valid~2 (
	.dataa(!out_data_4),
	.datab(!Equal16),
	.datac(!Equal14),
	.datad(!write_addr_data_both_valid),
	.datae(!src2_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src2_valid2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src2_valid~2 .extended_lut = "off";
defparam \src2_valid~2 .lut_mask = 64'h0002000000020000;
defparam \src2_valid~2 .shared_arith = "off";

cyclonev_lcell_comb \src6_valid~0 (
	.dataa(!has_pending_responses),
	.datab(!last_channel_6),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src6_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src6_valid~0 .extended_lut = "off";
defparam \src6_valid~0 .lut_mask = 64'h4444444444444444;
defparam \src6_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src6_valid~1 (
	.dataa(!write_addr_data_both_valid),
	.datab(!src6_valid),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src6_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src6_valid~1 .extended_lut = "off";
defparam \src6_valid~1 .lut_mask = 64'h4444444444444444;
defparam \src6_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \src6_valid~2 (
	.dataa(!out_data_4),
	.datab(!Equal5),
	.datac(!Equal14),
	.datad(!write_addr_data_both_valid),
	.datae(!src6_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src6_valid2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src6_valid~2 .extended_lut = "off";
defparam \src6_valid~2 .lut_mask = 64'h0002000000020000;
defparam \src6_valid~2 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~0 (
	.dataa(!out_data_5),
	.datab(!Equal15),
	.datac(!Equal13),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~0 .extended_lut = "off";
defparam \sink_ready~0 .lut_mask = 64'h0001000100010001;
defparam \sink_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~1 (
	.dataa(!out_data_4),
	.datab(!Equal16),
	.datac(!Equal161),
	.datad(!saved_grant_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_ready~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~1 .extended_lut = "off";
defparam \sink_ready~1 .lut_mask = 64'h0002000200020002;
defparam \sink_ready~1 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~2 (
	.dataa(!out_data_5),
	.datab(!Equal15),
	.datac(!Equal13),
	.datad(!saved_grant_02),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_ready~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~2 .extended_lut = "off";
defparam \sink_ready~2 .lut_mask = 64'h0002000200020002;
defparam \sink_ready~2 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~3 (
	.dataa(!out_data_4),
	.datab(!Equal14),
	.datac(!Equal13),
	.datad(!saved_grant_03),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_ready~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~3 .extended_lut = "off";
defparam \sink_ready~3 .lut_mask = 64'h0002000200020002;
defparam \sink_ready~3 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~4 (
	.dataa(!out_data_4),
	.datab(!Equal5),
	.datac(!Equal14),
	.datad(!saved_grant_04),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_ready~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~4 .extended_lut = "off";
defparam \sink_ready~4 .lut_mask = 64'h0002000200020002;
defparam \sink_ready~4 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~5 (
	.dataa(!out_data_5),
	.datab(!Equal15),
	.datac(!Equal9),
	.datad(!saved_grant_05),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_ready~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~5 .extended_lut = "off";
defparam \sink_ready~5 .lut_mask = 64'h0002000200020002;
defparam \sink_ready~5 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~6 (
	.dataa(!saved_grant_06),
	.datab(!out_data_8),
	.datac(!out_data_5),
	.datad(!out_data_4),
	.datae(!out_data_7),
	.dataf(!out_data_6),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_ready~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~6 .extended_lut = "off";
defparam \sink_ready~6 .lut_mask = 64'h4115551551155111;
defparam \sink_ready~6 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~7 (
	.dataa(!out_data_5),
	.datab(!Equal16),
	.datac(!Equal15),
	.datad(!saved_grant_07),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_ready~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~7 .extended_lut = "off";
defparam \sink_ready~7 .lut_mask = 64'h0002000200020002;
defparam \sink_ready~7 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~8 (
	.dataa(!out_data_4),
	.datab(!Equal16),
	.datac(!Equal14),
	.datad(!saved_grant_08),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_ready~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~8 .extended_lut = "off";
defparam \sink_ready~8 .lut_mask = 64'h0002000200020002;
defparam \sink_ready~8 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~9 (
	.dataa(!out_data_5),
	.datab(!Equal15),
	.datac(!Equal5),
	.datad(!saved_grant_09),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_ready~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~9 .extended_lut = "off";
defparam \sink_ready~9 .lut_mask = 64'h0002000200020002;
defparam \sink_ready~9 .shared_arith = "off";

cyclonev_lcell_comb \src0_valid~0 (
	.dataa(!h2f_AWVALID_0),
	.datab(!h2f_WVALID_0),
	.datac(!has_pending_responses),
	.datad(!last_channel_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src0_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src0_valid~0 .extended_lut = "off";
defparam \src0_valid~0 .lut_mask = 64'h1011101110111011;
defparam \src0_valid~0 .shared_arith = "off";

endmodule

module spw_babasu_spw_babasu_mm_interconnect_0_cmd_demux_1 (
	h2f_ARVALID_0,
	h2f_ARADDR_4,
	h2f_ARADDR_5,
	h2f_ARADDR_6,
	h2f_ARADDR_7,
	h2f_ARADDR_8,
	nxt_in_ready,
	nxt_in_ready1,
	nxt_in_ready2,
	nxt_in_ready3,
	nxt_in_ready4,
	nxt_in_ready5,
	nxt_in_ready6,
	nxt_in_ready7,
	nxt_in_ready8,
	nxt_in_ready9,
	has_pending_responses,
	last_channel_6,
	Equal6,
	saved_grant_1,
	stateST_COMP_TRANS,
	cp_ready,
	nxt_out_eop,
	src_channel,
	nxt_in_ready10,
	saved_grant_11,
	stateST_COMP_TRANS1,
	cp_ready1,
	nxt_out_eop1,
	last_cycle,
	nxt_in_ready11,
	saved_grant_12,
	stateST_COMP_TRANS2,
	cp_ready2,
	nxt_out_eop2,
	last_cycle1,
	nxt_in_ready12,
	nxt_in_ready13,
	saved_grant_13,
	src_channel_1,
	WideOr0,
	nxt_in_ready14,
	saved_grant_14,
	Equal15,
	nxt_in_ready15,
	Equal16,
	saved_grant_15,
	WideOr01,
	nxt_in_ready16,
	saved_grant_16,
	src_channel_13,
	nxt_in_ready17,
	saved_grant_17,
	Equal14,
	WideOr02,
	Equal3,
	saved_grant_18,
	stateST_COMP_TRANS3,
	cp_ready3,
	nxt_out_eop3,
	nxt_in_ready18,
	nxt_in_ready19,
	saved_grant_19,
	nxt_in_ready20,
	saved_grant_110,
	saved_grant_111,
	Equal10,
	stateST_COMP_TRANS4,
	cp_ready4,
	nxt_out_eop4,
	nxt_in_ready21,
	saved_grant_112,
	nxt_in_ready22,
	src_channel_0,
	nxt_in_ready23,
	nxt_in_ready24,
	nxt_in_ready25,
	saved_grant_113,
	nxt_in_ready26,
	saved_grant_114,
	nxt_in_ready27,
	saved_grant_115,
	nxt_in_ready28,
	saved_grant_116,
	WideOr03,
	last_channel_1,
	src1_valid,
	last_channel_15,
	src15_valid,
	src15_valid1,
	last_channel_16,
	src16_valid,
	src16_valid1,
	last_channel_14,
	src14_valid,
	src14_valid1,
	Equal9,
	last_channel_9,
	src9_valid,
	src9_valid1,
	last_channel_0,
	src0_valid,
	src_channel_2,
	last_channel_2,
	src2_valid,
	src2_valid1,
	src6_valid,
	src6_valid1)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARVALID_0;
input 	h2f_ARADDR_4;
input 	h2f_ARADDR_5;
input 	h2f_ARADDR_6;
input 	h2f_ARADDR_7;
input 	h2f_ARADDR_8;
input 	nxt_in_ready;
input 	nxt_in_ready1;
input 	nxt_in_ready2;
input 	nxt_in_ready3;
input 	nxt_in_ready4;
input 	nxt_in_ready5;
input 	nxt_in_ready6;
input 	nxt_in_ready7;
input 	nxt_in_ready8;
input 	nxt_in_ready9;
input 	has_pending_responses;
input 	last_channel_6;
input 	Equal6;
input 	saved_grant_1;
input 	stateST_COMP_TRANS;
input 	cp_ready;
input 	nxt_out_eop;
input 	src_channel;
input 	nxt_in_ready10;
input 	saved_grant_11;
input 	stateST_COMP_TRANS1;
input 	cp_ready1;
input 	nxt_out_eop1;
input 	last_cycle;
input 	nxt_in_ready11;
input 	saved_grant_12;
input 	stateST_COMP_TRANS2;
input 	cp_ready2;
input 	nxt_out_eop2;
input 	last_cycle1;
input 	nxt_in_ready12;
input 	nxt_in_ready13;
input 	saved_grant_13;
input 	src_channel_1;
output 	WideOr0;
input 	nxt_in_ready14;
input 	saved_grant_14;
input 	Equal15;
input 	nxt_in_ready15;
input 	Equal16;
input 	saved_grant_15;
output 	WideOr01;
input 	nxt_in_ready16;
input 	saved_grant_16;
input 	src_channel_13;
input 	nxt_in_ready17;
input 	saved_grant_17;
input 	Equal14;
output 	WideOr02;
input 	Equal3;
input 	saved_grant_18;
input 	stateST_COMP_TRANS3;
input 	cp_ready3;
input 	nxt_out_eop3;
input 	nxt_in_ready18;
input 	nxt_in_ready19;
input 	saved_grant_19;
input 	nxt_in_ready20;
input 	saved_grant_110;
input 	saved_grant_111;
input 	Equal10;
input 	stateST_COMP_TRANS4;
input 	cp_ready4;
input 	nxt_out_eop4;
input 	nxt_in_ready21;
input 	saved_grant_112;
input 	nxt_in_ready22;
input 	src_channel_0;
input 	nxt_in_ready23;
input 	nxt_in_ready24;
input 	nxt_in_ready25;
input 	saved_grant_113;
input 	nxt_in_ready26;
input 	saved_grant_114;
input 	nxt_in_ready27;
input 	saved_grant_115;
input 	nxt_in_ready28;
input 	saved_grant_116;
output 	WideOr03;
input 	last_channel_1;
output 	src1_valid;
input 	last_channel_15;
output 	src15_valid;
output 	src15_valid1;
input 	last_channel_16;
output 	src16_valid;
output 	src16_valid1;
input 	last_channel_14;
output 	src14_valid;
output 	src14_valid1;
input 	Equal9;
input 	last_channel_9;
output 	src9_valid;
output 	src9_valid1;
input 	last_channel_0;
output 	src0_valid;
input 	src_channel_2;
input 	last_channel_2;
output 	src2_valid;
output 	src2_valid1;
output 	src6_valid;
output 	src6_valid1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \sink_ready~0_combout ;
wire \sink_ready~1_combout ;
wire \sink_ready~2_combout ;
wire \sink_ready~3_combout ;
wire \sink_ready~4_combout ;
wire \sink_ready~5_combout ;
wire \sink_ready~6_combout ;
wire \sink_ready~7_combout ;
wire \sink_ready~8_combout ;
wire \sink_ready~9_combout ;
wire \sink_ready~10_combout ;
wire \WideOr0~3_combout ;
wire \sink_ready~11_combout ;
wire \sink_ready~12_combout ;
wire \sink_ready~13_combout ;
wire \sink_ready~14_combout ;
wire \WideOr0~4_combout ;
wire \sink_ready~15_combout ;
wire \sink_ready~16_combout ;
wire \WideOr0~5_combout ;


cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!\sink_ready~0_combout ),
	.datab(!\sink_ready~1_combout ),
	.datac(!\sink_ready~2_combout ),
	.datad(!nxt_in_ready13),
	.datae(!nxt_in_ready9),
	.dataf(!\sink_ready~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h8080808080000000;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~1 (
	.dataa(!nxt_in_ready14),
	.datab(!nxt_in_ready8),
	.datac(!\sink_ready~4_combout ),
	.datad(!nxt_in_ready15),
	.datae(!nxt_in_ready7),
	.dataf(!\sink_ready~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr01),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~1 .extended_lut = "off";
defparam \WideOr0~1 .lut_mask = 64'hF8F8F8F8F8000000;
defparam \WideOr0~1 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~2 (
	.dataa(!nxt_in_ready16),
	.datab(!nxt_in_ready6),
	.datac(!\sink_ready~6_combout ),
	.datad(!nxt_in_ready17),
	.datae(!nxt_in_ready5),
	.dataf(!\sink_ready~7_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr02),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~2 .extended_lut = "off";
defparam \WideOr0~2 .lut_mask = 64'hF8F8F8F8F8000000;
defparam \WideOr0~2 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~6 (
	.dataa(!\sink_ready~8_combout ),
	.datab(!\WideOr0~3_combout ),
	.datac(!\sink_ready~11_combout ),
	.datad(!\sink_ready~12_combout ),
	.datae(!\WideOr0~4_combout ),
	.dataf(!\WideOr0~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr03),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~6 .extended_lut = "off";
defparam \WideOr0~6 .lut_mask = 64'h0000000000002000;
defparam \WideOr0~6 .shared_arith = "off";

cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!h2f_ARVALID_0),
	.datab(!has_pending_responses),
	.datac(!src_channel_1),
	.datad(!last_channel_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'h0405040504050405;
defparam \src1_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src15_valid~0 (
	.dataa(!h2f_ARVALID_0),
	.datab(!has_pending_responses),
	.datac(!last_channel_15),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src15_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src15_valid~0 .extended_lut = "off";
defparam \src15_valid~0 .lut_mask = 64'h4545454545454545;
defparam \src15_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src15_valid~1 (
	.dataa(!Equal15),
	.datab(!src15_valid),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src15_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src15_valid~1 .extended_lut = "off";
defparam \src15_valid~1 .lut_mask = 64'h1111111111111111;
defparam \src15_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \src16_valid~0 (
	.dataa(!h2f_ARVALID_0),
	.datab(!has_pending_responses),
	.datac(!last_channel_16),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src16_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src16_valid~0 .extended_lut = "off";
defparam \src16_valid~0 .lut_mask = 64'h4545454545454545;
defparam \src16_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src16_valid~1 (
	.dataa(!Equal16),
	.datab(!src16_valid),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src16_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src16_valid~1 .extended_lut = "off";
defparam \src16_valid~1 .lut_mask = 64'h1111111111111111;
defparam \src16_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \src14_valid~0 (
	.dataa(!h2f_ARVALID_0),
	.datab(!has_pending_responses),
	.datac(!last_channel_14),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src14_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src14_valid~0 .extended_lut = "off";
defparam \src14_valid~0 .lut_mask = 64'h4545454545454545;
defparam \src14_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src14_valid~1 (
	.dataa(!Equal14),
	.datab(!src14_valid),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src14_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src14_valid~1 .extended_lut = "off";
defparam \src14_valid~1 .lut_mask = 64'h1111111111111111;
defparam \src14_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \src9_valid~0 (
	.dataa(!h2f_ARVALID_0),
	.datab(!has_pending_responses),
	.datac(!last_channel_9),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src9_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src9_valid~0 .extended_lut = "off";
defparam \src9_valid~0 .lut_mask = 64'h4545454545454545;
defparam \src9_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src9_valid~1 (
	.dataa(!Equal9),
	.datab(!src9_valid),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src9_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src9_valid~1 .extended_lut = "off";
defparam \src9_valid~1 .lut_mask = 64'h1111111111111111;
defparam \src9_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \src0_valid~0 (
	.dataa(!h2f_ARVALID_0),
	.datab(!has_pending_responses),
	.datac(!src_channel_0),
	.datad(!last_channel_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src0_valid~0 .extended_lut = "off";
defparam \src0_valid~0 .lut_mask = 64'h0405040504050405;
defparam \src0_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src2_valid~0 (
	.dataa(!h2f_ARVALID_0),
	.datab(!has_pending_responses),
	.datac(!last_channel_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src2_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src2_valid~0 .extended_lut = "off";
defparam \src2_valid~0 .lut_mask = 64'h4545454545454545;
defparam \src2_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src2_valid~1 (
	.dataa(!src_channel_2),
	.datab(!src2_valid),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src2_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src2_valid~1 .extended_lut = "off";
defparam \src2_valid~1 .lut_mask = 64'h1111111111111111;
defparam \src2_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \src6_valid~0 (
	.dataa(!h2f_ARVALID_0),
	.datab(!has_pending_responses),
	.datac(!last_channel_6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src6_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src6_valid~0 .extended_lut = "off";
defparam \src6_valid~0 .lut_mask = 64'h4545454545454545;
defparam \src6_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src6_valid~1 (
	.dataa(!Equal6),
	.datab(!src6_valid),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src6_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src6_valid~1 .extended_lut = "off";
defparam \src6_valid~1 .lut_mask = 64'h1111111111111111;
defparam \src6_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~0 (
	.dataa(!saved_grant_1),
	.datab(!stateST_COMP_TRANS),
	.datac(!cp_ready),
	.datad(!nxt_out_eop),
	.datae(!src_channel),
	.dataf(!nxt_in_ready10),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~0 .extended_lut = "off";
defparam \sink_ready~0 .lut_mask = 64'h0000555500000001;
defparam \sink_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~1 (
	.dataa(!saved_grant_11),
	.datab(!stateST_COMP_TRANS1),
	.datac(!cp_ready1),
	.datad(!nxt_out_eop1),
	.datae(!last_cycle),
	.dataf(!nxt_in_ready11),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_ready~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~1 .extended_lut = "off";
defparam \sink_ready~1 .lut_mask = 64'h0000555500000001;
defparam \sink_ready~1 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~2 (
	.dataa(!saved_grant_12),
	.datab(!stateST_COMP_TRANS2),
	.datac(!cp_ready2),
	.datad(!nxt_out_eop2),
	.datae(!last_cycle1),
	.dataf(!nxt_in_ready12),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_ready~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~2 .extended_lut = "off";
defparam \sink_ready~2 .lut_mask = 64'h0000555500000001;
defparam \sink_ready~2 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~3 (
	.dataa(!saved_grant_13),
	.datab(!src_channel_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_ready~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~3 .extended_lut = "off";
defparam \sink_ready~3 .lut_mask = 64'h1111111111111111;
defparam \sink_ready~3 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~4 (
	.dataa(!saved_grant_14),
	.datab(!Equal15),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_ready~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~4 .extended_lut = "off";
defparam \sink_ready~4 .lut_mask = 64'h1111111111111111;
defparam \sink_ready~4 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~5 (
	.dataa(!Equal16),
	.datab(!saved_grant_15),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_ready~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~5 .extended_lut = "off";
defparam \sink_ready~5 .lut_mask = 64'h1111111111111111;
defparam \sink_ready~5 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~6 (
	.dataa(!saved_grant_16),
	.datab(!src_channel_13),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_ready~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~6 .extended_lut = "off";
defparam \sink_ready~6 .lut_mask = 64'h1111111111111111;
defparam \sink_ready~6 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~7 (
	.dataa(!saved_grant_17),
	.datab(!Equal14),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_ready~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~7 .extended_lut = "off";
defparam \sink_ready~7 .lut_mask = 64'h1111111111111111;
defparam \sink_ready~7 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~8 (
	.dataa(!Equal3),
	.datab(!saved_grant_18),
	.datac(!stateST_COMP_TRANS3),
	.datad(!cp_ready3),
	.datae(!nxt_out_eop3),
	.dataf(!nxt_in_ready18),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_ready~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~8 .extended_lut = "off";
defparam \sink_ready~8 .lut_mask = 64'h1111111100000001;
defparam \sink_ready~8 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~9 (
	.dataa(!h2f_ARADDR_4),
	.datab(!h2f_ARADDR_5),
	.datac(!h2f_ARADDR_6),
	.datad(!h2f_ARADDR_7),
	.datae(!h2f_ARADDR_8),
	.dataf(!saved_grant_19),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_ready~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~9 .extended_lut = "off";
defparam \sink_ready~9 .lut_mask = 64'h0000000004000000;
defparam \sink_ready~9 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~10 (
	.dataa(!h2f_ARADDR_4),
	.datab(!h2f_ARADDR_5),
	.datac(!h2f_ARADDR_6),
	.datad(!h2f_ARADDR_7),
	.datae(!h2f_ARADDR_8),
	.dataf(!saved_grant_110),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_ready~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~10 .extended_lut = "off";
defparam \sink_ready~10 .lut_mask = 64'h0000000000400000;
defparam \sink_ready~10 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~3 (
	.dataa(!nxt_in_ready19),
	.datab(!nxt_in_ready4),
	.datac(!\sink_ready~9_combout ),
	.datad(!nxt_in_ready20),
	.datae(!nxt_in_ready3),
	.dataf(!\sink_ready~10_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~3 .extended_lut = "off";
defparam \WideOr0~3 .lut_mask = 64'hF8F8F8F8F8000000;
defparam \WideOr0~3 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~11 (
	.dataa(!saved_grant_111),
	.datab(!Equal10),
	.datac(!stateST_COMP_TRANS4),
	.datad(!cp_ready4),
	.datae(!nxt_out_eop4),
	.dataf(!nxt_in_ready21),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_ready~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~11 .extended_lut = "off";
defparam \sink_ready~11 .lut_mask = 64'h1111111100000001;
defparam \sink_ready~11 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~12 (
	.dataa(!saved_grant_112),
	.datab(!nxt_in_ready22),
	.datac(!nxt_in_ready2),
	.datad(!src_channel_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_ready~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~12 .extended_lut = "off";
defparam \sink_ready~12 .lut_mask = 64'h0015001500150015;
defparam \sink_ready~12 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~13 (
	.dataa(!h2f_ARADDR_4),
	.datab(!h2f_ARADDR_5),
	.datac(!h2f_ARADDR_6),
	.datad(!h2f_ARADDR_7),
	.datae(!h2f_ARADDR_8),
	.dataf(!saved_grant_113),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_ready~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~13 .extended_lut = "off";
defparam \sink_ready~13 .lut_mask = 64'h0000000008000000;
defparam \sink_ready~13 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~14 (
	.dataa(!h2f_ARADDR_4),
	.datab(!h2f_ARADDR_5),
	.datac(!h2f_ARADDR_6),
	.datad(!h2f_ARADDR_7),
	.datae(!h2f_ARADDR_8),
	.dataf(!saved_grant_114),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_ready~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~14 .extended_lut = "off";
defparam \sink_ready~14 .lut_mask = 64'h0000000001000000;
defparam \sink_ready~14 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~4 (
	.dataa(!nxt_in_ready23),
	.datab(!nxt_in_ready24),
	.datac(!nxt_in_ready25),
	.datad(!\sink_ready~13_combout ),
	.datae(!nxt_in_ready26),
	.dataf(!\sink_ready~14_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~4 .extended_lut = "off";
defparam \WideOr0~4 .lut_mask = 64'hFF0AFF0A0000CC08;
defparam \WideOr0~4 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~15 (
	.dataa(!h2f_ARADDR_4),
	.datab(!h2f_ARADDR_5),
	.datac(!h2f_ARADDR_6),
	.datad(!h2f_ARADDR_7),
	.datae(!h2f_ARADDR_8),
	.dataf(!saved_grant_115),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_ready~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~15 .extended_lut = "off";
defparam \sink_ready~15 .lut_mask = 64'h0000000020000000;
defparam \sink_ready~15 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~16 (
	.dataa(!h2f_ARADDR_4),
	.datab(!h2f_ARADDR_5),
	.datac(!h2f_ARADDR_6),
	.datad(!h2f_ARADDR_7),
	.datae(!h2f_ARADDR_8),
	.dataf(!saved_grant_116),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_ready~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~16 .extended_lut = "off";
defparam \sink_ready~16 .lut_mask = 64'h0000000002000000;
defparam \sink_ready~16 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~5 (
	.dataa(!nxt_in_ready27),
	.datab(!nxt_in_ready1),
	.datac(!\sink_ready~15_combout ),
	.datad(!nxt_in_ready28),
	.datae(!nxt_in_ready),
	.dataf(!\sink_ready~16_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~5 .extended_lut = "off";
defparam \WideOr0~5 .lut_mask = 64'hF8F8F8F8F8000000;
defparam \WideOr0~5 .shared_arith = "off";

endmodule

module spw_babasu_spw_babasu_mm_interconnect_0_cmd_mux (
	h2f_WLAST_0,
	h2f_ARID_0,
	h2f_ARID_1,
	h2f_ARID_2,
	h2f_ARID_3,
	h2f_ARID_4,
	h2f_ARID_5,
	h2f_ARID_6,
	h2f_ARID_7,
	h2f_ARID_8,
	h2f_ARID_9,
	h2f_ARID_10,
	h2f_ARID_11,
	h2f_ARSIZE_0,
	h2f_ARSIZE_1,
	h2f_ARSIZE_2,
	h2f_AWID_0,
	h2f_AWID_1,
	h2f_AWID_2,
	h2f_AWID_3,
	h2f_AWID_4,
	h2f_AWID_5,
	h2f_AWID_6,
	h2f_AWID_7,
	h2f_AWID_8,
	h2f_AWID_9,
	h2f_AWID_10,
	h2f_AWID_11,
	h2f_AWSIZE_0,
	h2f_AWSIZE_1,
	h2f_AWSIZE_2,
	h2f_WDATA_0,
	h2f_WSTRB_0,
	h2f_WSTRB_1,
	h2f_WSTRB_2,
	h2f_WSTRB_3,
	nxt_in_ready,
	saved_grant_1,
	nxt_in_ready1,
	saved_grant_0,
	altera_reset_synchronizer_int_chain_out,
	src0_valid,
	src0_valid1,
	nxt_in_ready2,
	src_valid,
	src_payload_0,
	src_data_87,
	src_data_88,
	src_data_35,
	src_data_34,
	src_data_33,
	src_data_32,
	Selector3,
	Selector10,
	Selector4,
	Selector11,
	src_payload,
	src_data_82,
	src_data_81,
	src_data_105,
	src_data_106,
	src_data_107,
	src_data_108,
	src_data_109,
	src_data_110,
	src_data_111,
	src_data_112,
	src_data_113,
	src_data_114,
	src_data_115,
	src_data_116,
	src_data_86,
	Selector5,
	Selector12,
	src_data_80,
	Selector6,
	Selector13,
	src_data_79,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_WLAST_0;
input 	h2f_ARID_0;
input 	h2f_ARID_1;
input 	h2f_ARID_2;
input 	h2f_ARID_3;
input 	h2f_ARID_4;
input 	h2f_ARID_5;
input 	h2f_ARID_6;
input 	h2f_ARID_7;
input 	h2f_ARID_8;
input 	h2f_ARID_9;
input 	h2f_ARID_10;
input 	h2f_ARID_11;
input 	h2f_ARSIZE_0;
input 	h2f_ARSIZE_1;
input 	h2f_ARSIZE_2;
input 	h2f_AWID_0;
input 	h2f_AWID_1;
input 	h2f_AWID_2;
input 	h2f_AWID_3;
input 	h2f_AWID_4;
input 	h2f_AWID_5;
input 	h2f_AWID_6;
input 	h2f_AWID_7;
input 	h2f_AWID_8;
input 	h2f_AWID_9;
input 	h2f_AWID_10;
input 	h2f_AWID_11;
input 	h2f_AWSIZE_0;
input 	h2f_AWSIZE_1;
input 	h2f_AWSIZE_2;
input 	h2f_WDATA_0;
input 	h2f_WSTRB_0;
input 	h2f_WSTRB_1;
input 	h2f_WSTRB_2;
input 	h2f_WSTRB_3;
input 	nxt_in_ready;
output 	saved_grant_1;
input 	nxt_in_ready1;
output 	saved_grant_0;
input 	altera_reset_synchronizer_int_chain_out;
input 	src0_valid;
input 	src0_valid1;
input 	nxt_in_ready2;
output 	src_valid;
output 	src_payload_0;
output 	src_data_87;
output 	src_data_88;
output 	src_data_35;
output 	src_data_34;
output 	src_data_33;
output 	src_data_32;
input 	Selector3;
input 	Selector10;
input 	Selector4;
input 	Selector11;
output 	src_payload;
output 	src_data_82;
output 	src_data_81;
output 	src_data_105;
output 	src_data_106;
output 	src_data_107;
output 	src_data_108;
output 	src_data_109;
output 	src_data_110;
output 	src_data_111;
output 	src_data_112;
output 	src_data_113;
output 	src_data_114;
output 	src_data_115;
output 	src_data_116;
output 	src_data_86;
input 	Selector5;
input 	Selector12;
output 	src_data_80;
input 	Selector6;
input 	Selector13;
output 	src_data_79;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[1]~0_combout ;
wire \arb|grant[0]~1_combout ;
wire \WideOr1~combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~0_combout ;


spw_babasu_altera_merlin_arbitrator_16 arb(
	.nxt_in_ready(nxt_in_ready),
	.nxt_in_ready1(nxt_in_ready1),
	.reset(altera_reset_synchronizer_int_chain_out),
	.src0_valid(src0_valid),
	.src0_valid1(src0_valid1),
	.grant_1(\arb|grant[1]~0_combout ),
	.src_payload_0(src_payload_0),
	.packet_in_progress(\packet_in_progress~q ),
	.grant_0(\arb|grant[0]~1_combout ),
	.WideOr1(\WideOr1~combout ),
	.clk(clk_clk));

cyclonev_lcell_comb WideOr1(
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!src0_valid),
	.datad(!src0_valid1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr1.extended_lut = "off";
defparam WideOr1.lut_mask = 64'h0357035703570357;
defparam WideOr1.shared_arith = "off";

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

cyclonev_lcell_comb \src_valid~0 (
	.dataa(!saved_grant_1),
	.datab(!src0_valid1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~0 .extended_lut = "off";
defparam \src_valid~0 .lut_mask = 64'h1111111111111111;
defparam \src_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload[0] (
	.dataa(!h2f_WLAST_0),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload[0] .extended_lut = "off";
defparam \src_payload[0] .lut_mask = 64'h3737373737373737;
defparam \src_payload[0] .shared_arith = "off";

cyclonev_lcell_comb \src_data[87] (
	.dataa(!h2f_ARSIZE_1),
	.datab(!h2f_AWSIZE_1),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_87),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[87] .extended_lut = "off";
defparam \src_data[87] .lut_mask = 64'h0537053705370537;
defparam \src_data[87] .shared_arith = "off";

cyclonev_lcell_comb \src_data[88] (
	.dataa(!h2f_ARSIZE_2),
	.datab(!h2f_AWSIZE_2),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_88),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[88] .extended_lut = "off";
defparam \src_data[88] .lut_mask = 64'h0537053705370537;
defparam \src_data[88] .shared_arith = "off";

cyclonev_lcell_comb \src_data[35] (
	.dataa(!h2f_WSTRB_3),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_35),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[35] .extended_lut = "off";
defparam \src_data[35] .lut_mask = 64'h3737373737373737;
defparam \src_data[35] .shared_arith = "off";

cyclonev_lcell_comb \src_data[34] (
	.dataa(!h2f_WSTRB_2),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_34),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[34] .extended_lut = "off";
defparam \src_data[34] .lut_mask = 64'h3737373737373737;
defparam \src_data[34] .shared_arith = "off";

cyclonev_lcell_comb \src_data[33] (
	.dataa(!h2f_WSTRB_1),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_33),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[33] .extended_lut = "off";
defparam \src_data[33] .lut_mask = 64'h3737373737373737;
defparam \src_data[33] .shared_arith = "off";

cyclonev_lcell_comb \src_data[32] (
	.dataa(!h2f_WSTRB_0),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_32),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[32] .extended_lut = "off";
defparam \src_data[32] .lut_mask = 64'h3737373737373737;
defparam \src_data[32] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!h2f_WDATA_0),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h1111111111111111;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[82] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector3),
	.datad(!Selector10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_82),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[82] .extended_lut = "off";
defparam \src_data[82] .lut_mask = 64'h0357035703570357;
defparam \src_data[82] .shared_arith = "off";

cyclonev_lcell_comb \src_data[81] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector4),
	.datad(!Selector11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_81),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[81] .extended_lut = "off";
defparam \src_data[81] .lut_mask = 64'h0357035703570357;
defparam \src_data[81] .shared_arith = "off";

cyclonev_lcell_comb \src_data[105] (
	.dataa(!h2f_ARID_0),
	.datab(!h2f_AWID_0),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_105),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[105] .extended_lut = "off";
defparam \src_data[105] .lut_mask = 64'h0537053705370537;
defparam \src_data[105] .shared_arith = "off";

cyclonev_lcell_comb \src_data[106] (
	.dataa(!h2f_ARID_1),
	.datab(!h2f_AWID_1),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_106),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[106] .extended_lut = "off";
defparam \src_data[106] .lut_mask = 64'h0537053705370537;
defparam \src_data[106] .shared_arith = "off";

cyclonev_lcell_comb \src_data[107] (
	.dataa(!h2f_ARID_2),
	.datab(!h2f_AWID_2),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_107),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[107] .extended_lut = "off";
defparam \src_data[107] .lut_mask = 64'h0537053705370537;
defparam \src_data[107] .shared_arith = "off";

cyclonev_lcell_comb \src_data[108] (
	.dataa(!h2f_ARID_3),
	.datab(!h2f_AWID_3),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_108),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[108] .extended_lut = "off";
defparam \src_data[108] .lut_mask = 64'h0537053705370537;
defparam \src_data[108] .shared_arith = "off";

cyclonev_lcell_comb \src_data[109] (
	.dataa(!h2f_ARID_4),
	.datab(!h2f_AWID_4),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_109),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[109] .extended_lut = "off";
defparam \src_data[109] .lut_mask = 64'h0537053705370537;
defparam \src_data[109] .shared_arith = "off";

cyclonev_lcell_comb \src_data[110] (
	.dataa(!h2f_ARID_5),
	.datab(!h2f_AWID_5),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_110),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[110] .extended_lut = "off";
defparam \src_data[110] .lut_mask = 64'h0537053705370537;
defparam \src_data[110] .shared_arith = "off";

cyclonev_lcell_comb \src_data[111] (
	.dataa(!h2f_ARID_6),
	.datab(!h2f_AWID_6),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_111),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[111] .extended_lut = "off";
defparam \src_data[111] .lut_mask = 64'h0537053705370537;
defparam \src_data[111] .shared_arith = "off";

cyclonev_lcell_comb \src_data[112] (
	.dataa(!h2f_ARID_7),
	.datab(!h2f_AWID_7),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_112),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[112] .extended_lut = "off";
defparam \src_data[112] .lut_mask = 64'h0537053705370537;
defparam \src_data[112] .shared_arith = "off";

cyclonev_lcell_comb \src_data[113] (
	.dataa(!h2f_ARID_8),
	.datab(!h2f_AWID_8),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_113),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[113] .extended_lut = "off";
defparam \src_data[113] .lut_mask = 64'h0537053705370537;
defparam \src_data[113] .shared_arith = "off";

cyclonev_lcell_comb \src_data[114] (
	.dataa(!h2f_ARID_9),
	.datab(!h2f_AWID_9),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_114),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[114] .extended_lut = "off";
defparam \src_data[114] .lut_mask = 64'h0537053705370537;
defparam \src_data[114] .shared_arith = "off";

cyclonev_lcell_comb \src_data[115] (
	.dataa(!h2f_ARID_10),
	.datab(!h2f_AWID_10),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_115),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[115] .extended_lut = "off";
defparam \src_data[115] .lut_mask = 64'h0537053705370537;
defparam \src_data[115] .shared_arith = "off";

cyclonev_lcell_comb \src_data[116] (
	.dataa(!h2f_ARID_11),
	.datab(!h2f_AWID_11),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_116),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[116] .extended_lut = "off";
defparam \src_data[116] .lut_mask = 64'h0537053705370537;
defparam \src_data[116] .shared_arith = "off";

cyclonev_lcell_comb \src_data[86] (
	.dataa(!h2f_ARSIZE_0),
	.datab(!h2f_AWSIZE_0),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_86),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[86] .extended_lut = "off";
defparam \src_data[86] .lut_mask = 64'h0537053705370537;
defparam \src_data[86] .shared_arith = "off";

cyclonev_lcell_comb \src_data[80] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector5),
	.datad(!Selector12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_80),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[80] .extended_lut = "off";
defparam \src_data[80] .lut_mask = 64'h0357035703570357;
defparam \src_data[80] .shared_arith = "off";

cyclonev_lcell_comb \src_data[79] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector6),
	.datad(!Selector13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_79),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[79] .extended_lut = "off";
defparam \src_data[79] .lut_mask = 64'h0357035703570357;
defparam \src_data[79] .shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!\update_grant~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \update_grant~0 (
	.dataa(!nxt_in_ready2),
	.datab(!saved_grant_0),
	.datac(!src0_valid),
	.datad(!src_valid),
	.datae(!src_payload_0),
	.dataf(!\packet_in_progress~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\update_grant~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \update_grant~0 .extended_lut = "off";
defparam \update_grant~0 .lut_mask = 64'hFC00FEAA000002AA;
defparam \update_grant~0 .shared_arith = "off";

endmodule

module spw_babasu_spw_babasu_mm_interconnect_0_cmd_mux_1 (
	h2f_ARVALID_0,
	h2f_WLAST_0,
	h2f_ARID_0,
	h2f_ARID_1,
	h2f_ARID_2,
	h2f_ARID_3,
	h2f_ARID_4,
	h2f_ARID_5,
	h2f_ARID_6,
	h2f_ARID_7,
	h2f_ARID_8,
	h2f_ARID_9,
	h2f_ARID_10,
	h2f_ARID_11,
	h2f_ARSIZE_0,
	h2f_ARSIZE_1,
	h2f_ARSIZE_2,
	h2f_AWID_0,
	h2f_AWID_1,
	h2f_AWID_2,
	h2f_AWID_3,
	h2f_AWID_4,
	h2f_AWID_5,
	h2f_AWID_6,
	h2f_AWID_7,
	h2f_AWID_8,
	h2f_AWID_9,
	h2f_AWID_10,
	h2f_AWID_11,
	h2f_AWSIZE_0,
	h2f_AWSIZE_1,
	h2f_AWSIZE_2,
	h2f_WDATA_0,
	h2f_WSTRB_0,
	h2f_WSTRB_1,
	h2f_WSTRB_2,
	h2f_WSTRB_3,
	nxt_in_ready,
	has_pending_responses,
	nxt_in_ready1,
	saved_grant_1,
	src_channel_1,
	write_addr_data_both_valid,
	out_data_5,
	Equal16,
	Equal15,
	saved_grant_0,
	altera_reset_synchronizer_int_chain_out,
	Equal5,
	src1_valid,
	src1_valid1,
	last_channel_1,
	src_valid,
	src_data_87,
	src_data_88,
	src_valid1,
	src_data_35,
	src_data_34,
	src_data_33,
	src_data_32,
	src_payload_0,
	src1_valid2,
	src1_valid3,
	Selector3,
	Selector10,
	Selector4,
	Selector11,
	src_payload,
	src_data_82,
	src_data_81,
	src_data_105,
	src_data_106,
	src_data_107,
	src_data_108,
	src_data_109,
	src_data_110,
	src_data_111,
	src_data_112,
	src_data_113,
	src_data_114,
	src_data_115,
	src_data_116,
	src_data_86,
	Selector5,
	Selector12,
	src_data_80,
	Selector6,
	Selector13,
	src_data_79,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARVALID_0;
input 	h2f_WLAST_0;
input 	h2f_ARID_0;
input 	h2f_ARID_1;
input 	h2f_ARID_2;
input 	h2f_ARID_3;
input 	h2f_ARID_4;
input 	h2f_ARID_5;
input 	h2f_ARID_6;
input 	h2f_ARID_7;
input 	h2f_ARID_8;
input 	h2f_ARID_9;
input 	h2f_ARID_10;
input 	h2f_ARID_11;
input 	h2f_ARSIZE_0;
input 	h2f_ARSIZE_1;
input 	h2f_ARSIZE_2;
input 	h2f_AWID_0;
input 	h2f_AWID_1;
input 	h2f_AWID_2;
input 	h2f_AWID_3;
input 	h2f_AWID_4;
input 	h2f_AWID_5;
input 	h2f_AWID_6;
input 	h2f_AWID_7;
input 	h2f_AWID_8;
input 	h2f_AWID_9;
input 	h2f_AWID_10;
input 	h2f_AWID_11;
input 	h2f_AWSIZE_0;
input 	h2f_AWSIZE_1;
input 	h2f_AWSIZE_2;
input 	h2f_WDATA_0;
input 	h2f_WSTRB_0;
input 	h2f_WSTRB_1;
input 	h2f_WSTRB_2;
input 	h2f_WSTRB_3;
input 	nxt_in_ready;
input 	has_pending_responses;
input 	nxt_in_ready1;
output 	saved_grant_1;
input 	src_channel_1;
input 	write_addr_data_both_valid;
input 	out_data_5;
input 	Equal16;
input 	Equal15;
output 	saved_grant_0;
input 	altera_reset_synchronizer_int_chain_out;
input 	Equal5;
input 	src1_valid;
input 	src1_valid1;
input 	last_channel_1;
output 	src_valid;
output 	src_data_87;
output 	src_data_88;
output 	src_valid1;
output 	src_data_35;
output 	src_data_34;
output 	src_data_33;
output 	src_data_32;
output 	src_payload_0;
input 	src1_valid2;
input 	src1_valid3;
input 	Selector3;
input 	Selector10;
input 	Selector4;
input 	Selector11;
output 	src_payload;
output 	src_data_82;
output 	src_data_81;
output 	src_data_105;
output 	src_data_106;
output 	src_data_107;
output 	src_data_108;
output 	src_data_109;
output 	src_data_110;
output 	src_data_111;
output 	src_data_112;
output 	src_data_113;
output 	src_data_114;
output 	src_data_115;
output 	src_data_116;
output 	src_data_86;
input 	Selector5;
input 	Selector12;
output 	src_data_80;
input 	Selector6;
input 	Selector13;
output 	src_data_79;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[1]~0_combout ;
wire \arb|grant[0]~1_combout ;
wire \WideOr1~combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~0_combout ;


spw_babasu_altera_merlin_arbitrator arb(
	.nxt_in_ready(nxt_in_ready),
	.nxt_in_ready1(nxt_in_ready1),
	.write_addr_data_both_valid(write_addr_data_both_valid),
	.out_data_5(out_data_5),
	.Equal16(Equal16),
	.Equal15(Equal15),
	.reset(altera_reset_synchronizer_int_chain_out),
	.src1_valid(src1_valid),
	.src_payload_0(src_payload_0),
	.src1_valid1(src1_valid2),
	.src1_valid2(src1_valid3),
	.grant_1(\arb|grant[1]~0_combout ),
	.packet_in_progress(\packet_in_progress~q ),
	.grant_0(\arb|grant[0]~1_combout ),
	.WideOr1(\WideOr1~combout ),
	.clk(clk_clk));

cyclonev_lcell_comb WideOr1(
	.dataa(!Equal16),
	.datab(!Equal5),
	.datac(!saved_grant_0),
	.datad(!src1_valid1),
	.datae(!src_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr1.extended_lut = "off";
defparam WideOr1.lut_mask = 64'hFFFE0000FFFE0000;
defparam WideOr1.shared_arith = "off";

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

cyclonev_lcell_comb \src_valid~0 (
	.dataa(!h2f_ARVALID_0),
	.datab(!has_pending_responses),
	.datac(!saved_grant_1),
	.datad(!src_channel_1),
	.datae(!last_channel_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~0 .extended_lut = "off";
defparam \src_valid~0 .lut_mask = 64'h0004000500040005;
defparam \src_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[87] (
	.dataa(!h2f_ARSIZE_1),
	.datab(!h2f_AWSIZE_1),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_87),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[87] .extended_lut = "off";
defparam \src_data[87] .lut_mask = 64'h0537053705370537;
defparam \src_data[87] .shared_arith = "off";

cyclonev_lcell_comb \src_data[88] (
	.dataa(!h2f_ARSIZE_2),
	.datab(!h2f_AWSIZE_2),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_88),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[88] .extended_lut = "off";
defparam \src_data[88] .lut_mask = 64'h0537053705370537;
defparam \src_data[88] .shared_arith = "off";

cyclonev_lcell_comb \src_valid~1 (
	.dataa(!out_data_5),
	.datab(!Equal16),
	.datac(!Equal15),
	.datad(!saved_grant_0),
	.datae(!write_addr_data_both_valid),
	.dataf(!src1_valid),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~1 .extended_lut = "off";
defparam \src_valid~1 .lut_mask = 64'h0000000200000000;
defparam \src_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \src_data[35] (
	.dataa(!h2f_WSTRB_3),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_35),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[35] .extended_lut = "off";
defparam \src_data[35] .lut_mask = 64'h3737373737373737;
defparam \src_data[35] .shared_arith = "off";

cyclonev_lcell_comb \src_data[34] (
	.dataa(!h2f_WSTRB_2),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_34),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[34] .extended_lut = "off";
defparam \src_data[34] .lut_mask = 64'h3737373737373737;
defparam \src_data[34] .shared_arith = "off";

cyclonev_lcell_comb \src_data[33] (
	.dataa(!h2f_WSTRB_1),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_33),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[33] .extended_lut = "off";
defparam \src_data[33] .lut_mask = 64'h3737373737373737;
defparam \src_data[33] .shared_arith = "off";

cyclonev_lcell_comb \src_data[32] (
	.dataa(!h2f_WSTRB_0),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_32),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[32] .extended_lut = "off";
defparam \src_data[32] .lut_mask = 64'h3737373737373737;
defparam \src_data[32] .shared_arith = "off";

cyclonev_lcell_comb \src_payload[0] (
	.dataa(!h2f_WLAST_0),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload[0] .extended_lut = "off";
defparam \src_payload[0] .lut_mask = 64'h3737373737373737;
defparam \src_payload[0] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!h2f_WDATA_0),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h1111111111111111;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[82] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector3),
	.datad(!Selector10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_82),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[82] .extended_lut = "off";
defparam \src_data[82] .lut_mask = 64'h0357035703570357;
defparam \src_data[82] .shared_arith = "off";

cyclonev_lcell_comb \src_data[81] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector4),
	.datad(!Selector11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_81),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[81] .extended_lut = "off";
defparam \src_data[81] .lut_mask = 64'h0357035703570357;
defparam \src_data[81] .shared_arith = "off";

cyclonev_lcell_comb \src_data[105] (
	.dataa(!h2f_ARID_0),
	.datab(!h2f_AWID_0),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_105),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[105] .extended_lut = "off";
defparam \src_data[105] .lut_mask = 64'h0537053705370537;
defparam \src_data[105] .shared_arith = "off";

cyclonev_lcell_comb \src_data[106] (
	.dataa(!h2f_ARID_1),
	.datab(!h2f_AWID_1),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_106),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[106] .extended_lut = "off";
defparam \src_data[106] .lut_mask = 64'h0537053705370537;
defparam \src_data[106] .shared_arith = "off";

cyclonev_lcell_comb \src_data[107] (
	.dataa(!h2f_ARID_2),
	.datab(!h2f_AWID_2),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_107),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[107] .extended_lut = "off";
defparam \src_data[107] .lut_mask = 64'h0537053705370537;
defparam \src_data[107] .shared_arith = "off";

cyclonev_lcell_comb \src_data[108] (
	.dataa(!h2f_ARID_3),
	.datab(!h2f_AWID_3),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_108),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[108] .extended_lut = "off";
defparam \src_data[108] .lut_mask = 64'h0537053705370537;
defparam \src_data[108] .shared_arith = "off";

cyclonev_lcell_comb \src_data[109] (
	.dataa(!h2f_ARID_4),
	.datab(!h2f_AWID_4),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_109),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[109] .extended_lut = "off";
defparam \src_data[109] .lut_mask = 64'h0537053705370537;
defparam \src_data[109] .shared_arith = "off";

cyclonev_lcell_comb \src_data[110] (
	.dataa(!h2f_ARID_5),
	.datab(!h2f_AWID_5),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_110),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[110] .extended_lut = "off";
defparam \src_data[110] .lut_mask = 64'h0537053705370537;
defparam \src_data[110] .shared_arith = "off";

cyclonev_lcell_comb \src_data[111] (
	.dataa(!h2f_ARID_6),
	.datab(!h2f_AWID_6),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_111),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[111] .extended_lut = "off";
defparam \src_data[111] .lut_mask = 64'h0537053705370537;
defparam \src_data[111] .shared_arith = "off";

cyclonev_lcell_comb \src_data[112] (
	.dataa(!h2f_ARID_7),
	.datab(!h2f_AWID_7),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_112),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[112] .extended_lut = "off";
defparam \src_data[112] .lut_mask = 64'h0537053705370537;
defparam \src_data[112] .shared_arith = "off";

cyclonev_lcell_comb \src_data[113] (
	.dataa(!h2f_ARID_8),
	.datab(!h2f_AWID_8),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_113),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[113] .extended_lut = "off";
defparam \src_data[113] .lut_mask = 64'h0537053705370537;
defparam \src_data[113] .shared_arith = "off";

cyclonev_lcell_comb \src_data[114] (
	.dataa(!h2f_ARID_9),
	.datab(!h2f_AWID_9),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_114),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[114] .extended_lut = "off";
defparam \src_data[114] .lut_mask = 64'h0537053705370537;
defparam \src_data[114] .shared_arith = "off";

cyclonev_lcell_comb \src_data[115] (
	.dataa(!h2f_ARID_10),
	.datab(!h2f_AWID_10),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_115),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[115] .extended_lut = "off";
defparam \src_data[115] .lut_mask = 64'h0537053705370537;
defparam \src_data[115] .shared_arith = "off";

cyclonev_lcell_comb \src_data[116] (
	.dataa(!h2f_ARID_11),
	.datab(!h2f_AWID_11),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_116),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[116] .extended_lut = "off";
defparam \src_data[116] .lut_mask = 64'h0537053705370537;
defparam \src_data[116] .shared_arith = "off";

cyclonev_lcell_comb \src_data[86] (
	.dataa(!h2f_ARSIZE_0),
	.datab(!h2f_AWSIZE_0),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_86),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[86] .extended_lut = "off";
defparam \src_data[86] .lut_mask = 64'h0537053705370537;
defparam \src_data[86] .shared_arith = "off";

cyclonev_lcell_comb \src_data[80] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector5),
	.datad(!Selector12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_80),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[80] .extended_lut = "off";
defparam \src_data[80] .lut_mask = 64'h0357035703570357;
defparam \src_data[80] .shared_arith = "off";

cyclonev_lcell_comb \src_data[79] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector6),
	.datad(!Selector13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_79),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[79] .extended_lut = "off";
defparam \src_data[79] .lut_mask = 64'h0357035703570357;
defparam \src_data[79] .shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!\update_grant~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \update_grant~0 (
	.dataa(!nxt_in_ready1),
	.datab(!nxt_in_ready),
	.datac(!src_valid),
	.datad(!src_valid1),
	.datae(!src_payload_0),
	.dataf(!\packet_in_progress~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\update_grant~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \update_grant~0 .extended_lut = "off";
defparam \update_grant~0 .lut_mask = 64'hF000F77700000777;
defparam \update_grant~0 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_arbitrator (
	nxt_in_ready,
	nxt_in_ready1,
	write_addr_data_both_valid,
	out_data_5,
	Equal16,
	Equal15,
	reset,
	src1_valid,
	src_payload_0,
	src1_valid1,
	src1_valid2,
	grant_1,
	packet_in_progress,
	grant_0,
	WideOr1,
	clk)/* synthesis synthesis_greybox=0 */;
input 	nxt_in_ready;
input 	nxt_in_ready1;
input 	write_addr_data_both_valid;
input 	out_data_5;
input 	Equal16;
input 	Equal15;
input 	reset;
input 	src1_valid;
input 	src_payload_0;
input 	src1_valid1;
input 	src1_valid2;
output 	grant_1;
input 	packet_in_progress;
output 	grant_0;
input 	WideOr1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg[0]~2_combout ;
wire \top_priority_reg[0]~q ;


cyclonev_lcell_comb \grant[1]~0 (
	.dataa(!\top_priority_reg[1]~q ),
	.datab(!\top_priority_reg[0]~q ),
	.datac(!src1_valid1),
	.datad(!src1_valid2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[1]~0 .extended_lut = "off";
defparam \grant[1]~0 .lut_mask = 64'h00D500D500D500D5;
defparam \grant[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \grant[0]~1 (
	.dataa(!\top_priority_reg[1]~q ),
	.datab(!\top_priority_reg[0]~q ),
	.datac(!src1_valid1),
	.datad(!src1_valid2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[0]~1 .extended_lut = "off";
defparam \grant[0]~1 .lut_mask = 64'h0D0C0D0C0D0C0D0C;
defparam \grant[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~0 (
	.dataa(!out_data_5),
	.datab(!Equal16),
	.datac(!Equal15),
	.datad(!write_addr_data_both_valid),
	.datae(!src1_valid),
	.dataf(!src1_valid2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~0 .extended_lut = "off";
defparam \top_priority_reg[0]~0 .lut_mask = 64'hFFFDFFFF00000000;
defparam \top_priority_reg[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~1 (
	.dataa(!nxt_in_ready1),
	.datab(!nxt_in_ready),
	.datac(!WideOr1),
	.datad(!src_payload_0),
	.datae(!packet_in_progress),
	.dataf(!\top_priority_reg[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~1 .extended_lut = "off";
defparam \top_priority_reg[0]~1 .lut_mask = 64'h0F7F007000000000;
defparam \top_priority_reg[0]~1 .shared_arith = "off";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~1_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

cyclonev_lcell_comb \top_priority_reg[0]~2 (
	.dataa(!grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~2 .extended_lut = "off";
defparam \top_priority_reg[0]~2 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \top_priority_reg[0]~2 .shared_arith = "off";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~1_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

endmodule

module spw_babasu_spw_babasu_mm_interconnect_0_cmd_mux_2 (
	h2f_WLAST_0,
	h2f_ARID_0,
	h2f_ARID_1,
	h2f_ARID_2,
	h2f_ARID_3,
	h2f_ARID_4,
	h2f_ARID_5,
	h2f_ARID_6,
	h2f_ARID_7,
	h2f_ARID_8,
	h2f_ARID_9,
	h2f_ARID_10,
	h2f_ARID_11,
	h2f_ARSIZE_0,
	h2f_ARSIZE_1,
	h2f_ARSIZE_2,
	h2f_AWID_0,
	h2f_AWID_1,
	h2f_AWID_2,
	h2f_AWID_3,
	h2f_AWID_4,
	h2f_AWID_5,
	h2f_AWID_6,
	h2f_AWID_7,
	h2f_AWID_8,
	h2f_AWID_9,
	h2f_AWID_10,
	h2f_AWID_11,
	h2f_AWSIZE_0,
	h2f_AWSIZE_1,
	h2f_AWSIZE_2,
	h2f_WDATA_0,
	h2f_WSTRB_0,
	h2f_WSTRB_1,
	h2f_WSTRB_2,
	h2f_WSTRB_3,
	nxt_in_ready,
	nxt_in_ready1,
	saved_grant_1,
	write_addr_data_both_valid,
	out_data_4,
	Equal14,
	Equal16,
	saved_grant_0,
	altera_reset_synchronizer_int_chain_out,
	Equal141,
	src2_valid,
	src2_valid1,
	src_channel_2,
	src2_valid2,
	src_valid,
	src_data_87,
	src_data_88,
	src_valid1,
	src_data_35,
	src_data_34,
	src_data_33,
	src_data_32,
	src_payload_0,
	src2_valid3,
	src2_valid4,
	src_payload,
	Selector3,
	Selector10,
	src_data_82,
	Selector4,
	Selector11,
	src_data_81,
	src_data_105,
	src_data_106,
	src_data_107,
	src_data_108,
	src_data_109,
	src_data_110,
	src_data_111,
	src_data_112,
	src_data_113,
	src_data_114,
	src_data_115,
	src_data_116,
	src_data_86,
	Selector5,
	Selector12,
	src_data_80,
	Selector6,
	Selector13,
	src_data_79,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_WLAST_0;
input 	h2f_ARID_0;
input 	h2f_ARID_1;
input 	h2f_ARID_2;
input 	h2f_ARID_3;
input 	h2f_ARID_4;
input 	h2f_ARID_5;
input 	h2f_ARID_6;
input 	h2f_ARID_7;
input 	h2f_ARID_8;
input 	h2f_ARID_9;
input 	h2f_ARID_10;
input 	h2f_ARID_11;
input 	h2f_ARSIZE_0;
input 	h2f_ARSIZE_1;
input 	h2f_ARSIZE_2;
input 	h2f_AWID_0;
input 	h2f_AWID_1;
input 	h2f_AWID_2;
input 	h2f_AWID_3;
input 	h2f_AWID_4;
input 	h2f_AWID_5;
input 	h2f_AWID_6;
input 	h2f_AWID_7;
input 	h2f_AWID_8;
input 	h2f_AWID_9;
input 	h2f_AWID_10;
input 	h2f_AWID_11;
input 	h2f_AWSIZE_0;
input 	h2f_AWSIZE_1;
input 	h2f_AWSIZE_2;
input 	h2f_WDATA_0;
input 	h2f_WSTRB_0;
input 	h2f_WSTRB_1;
input 	h2f_WSTRB_2;
input 	h2f_WSTRB_3;
input 	nxt_in_ready;
input 	nxt_in_ready1;
output 	saved_grant_1;
input 	write_addr_data_both_valid;
input 	out_data_4;
input 	Equal14;
input 	Equal16;
output 	saved_grant_0;
input 	altera_reset_synchronizer_int_chain_out;
input 	Equal141;
input 	src2_valid;
input 	src2_valid1;
input 	src_channel_2;
input 	src2_valid2;
output 	src_valid;
output 	src_data_87;
output 	src_data_88;
output 	src_valid1;
output 	src_data_35;
output 	src_data_34;
output 	src_data_33;
output 	src_data_32;
output 	src_payload_0;
input 	src2_valid3;
input 	src2_valid4;
output 	src_payload;
input 	Selector3;
input 	Selector10;
output 	src_data_82;
input 	Selector4;
input 	Selector11;
output 	src_data_81;
output 	src_data_105;
output 	src_data_106;
output 	src_data_107;
output 	src_data_108;
output 	src_data_109;
output 	src_data_110;
output 	src_data_111;
output 	src_data_112;
output 	src_data_113;
output 	src_data_114;
output 	src_data_115;
output 	src_data_116;
output 	src_data_86;
input 	Selector5;
input 	Selector12;
output 	src_data_80;
input 	Selector6;
input 	Selector13;
output 	src_data_79;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[1]~0_combout ;
wire \arb|grant[0]~1_combout ;
wire \WideOr1~combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~0_combout ;


spw_babasu_altera_merlin_arbitrator_1 arb(
	.nxt_in_ready(nxt_in_ready),
	.nxt_in_ready1(nxt_in_ready1),
	.Equal16(Equal16),
	.reset(altera_reset_synchronizer_int_chain_out),
	.Equal14(Equal141),
	.src2_valid(src2_valid1),
	.src_payload_0(src_payload_0),
	.src2_valid1(src2_valid3),
	.src2_valid2(src2_valid4),
	.grant_1(\arb|grant[1]~0_combout ),
	.packet_in_progress(\packet_in_progress~q ),
	.grant_0(\arb|grant[0]~1_combout ),
	.WideOr1(\WideOr1~combout ),
	.clk(clk_clk));

cyclonev_lcell_comb WideOr1(
	.dataa(!Equal16),
	.datab(!Equal141),
	.datac(!saved_grant_0),
	.datad(!src2_valid1),
	.datae(!src_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr1.extended_lut = "off";
defparam WideOr1.lut_mask = 64'hFFFE0000FFFE0000;
defparam WideOr1.shared_arith = "off";

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

cyclonev_lcell_comb \src_valid~0 (
	.dataa(!saved_grant_1),
	.datab(!src_channel_2),
	.datac(!src2_valid2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~0 .extended_lut = "off";
defparam \src_valid~0 .lut_mask = 64'h0101010101010101;
defparam \src_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[87] (
	.dataa(!h2f_ARSIZE_1),
	.datab(!h2f_AWSIZE_1),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_87),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[87] .extended_lut = "off";
defparam \src_data[87] .lut_mask = 64'h0537053705370537;
defparam \src_data[87] .shared_arith = "off";

cyclonev_lcell_comb \src_data[88] (
	.dataa(!h2f_ARSIZE_2),
	.datab(!h2f_AWSIZE_2),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_88),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[88] .extended_lut = "off";
defparam \src_data[88] .lut_mask = 64'h0537053705370537;
defparam \src_data[88] .shared_arith = "off";

cyclonev_lcell_comb \src_valid~1 (
	.dataa(!out_data_4),
	.datab(!Equal16),
	.datac(!Equal14),
	.datad(!saved_grant_0),
	.datae(!write_addr_data_both_valid),
	.dataf(!src2_valid),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~1 .extended_lut = "off";
defparam \src_valid~1 .lut_mask = 64'h0000000200000000;
defparam \src_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \src_data[35] (
	.dataa(!h2f_WSTRB_3),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_35),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[35] .extended_lut = "off";
defparam \src_data[35] .lut_mask = 64'h3737373737373737;
defparam \src_data[35] .shared_arith = "off";

cyclonev_lcell_comb \src_data[34] (
	.dataa(!h2f_WSTRB_2),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_34),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[34] .extended_lut = "off";
defparam \src_data[34] .lut_mask = 64'h3737373737373737;
defparam \src_data[34] .shared_arith = "off";

cyclonev_lcell_comb \src_data[33] (
	.dataa(!h2f_WSTRB_1),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_33),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[33] .extended_lut = "off";
defparam \src_data[33] .lut_mask = 64'h3737373737373737;
defparam \src_data[33] .shared_arith = "off";

cyclonev_lcell_comb \src_data[32] (
	.dataa(!h2f_WSTRB_0),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_32),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[32] .extended_lut = "off";
defparam \src_data[32] .lut_mask = 64'h3737373737373737;
defparam \src_data[32] .shared_arith = "off";

cyclonev_lcell_comb \src_payload[0] (
	.dataa(!h2f_WLAST_0),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload[0] .extended_lut = "off";
defparam \src_payload[0] .lut_mask = 64'h3737373737373737;
defparam \src_payload[0] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!h2f_WDATA_0),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h1111111111111111;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[82] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector3),
	.datad(!Selector10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_82),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[82] .extended_lut = "off";
defparam \src_data[82] .lut_mask = 64'h0357035703570357;
defparam \src_data[82] .shared_arith = "off";

cyclonev_lcell_comb \src_data[81] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector4),
	.datad(!Selector11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_81),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[81] .extended_lut = "off";
defparam \src_data[81] .lut_mask = 64'h0357035703570357;
defparam \src_data[81] .shared_arith = "off";

cyclonev_lcell_comb \src_data[105] (
	.dataa(!h2f_ARID_0),
	.datab(!h2f_AWID_0),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_105),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[105] .extended_lut = "off";
defparam \src_data[105] .lut_mask = 64'h0537053705370537;
defparam \src_data[105] .shared_arith = "off";

cyclonev_lcell_comb \src_data[106] (
	.dataa(!h2f_ARID_1),
	.datab(!h2f_AWID_1),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_106),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[106] .extended_lut = "off";
defparam \src_data[106] .lut_mask = 64'h0537053705370537;
defparam \src_data[106] .shared_arith = "off";

cyclonev_lcell_comb \src_data[107] (
	.dataa(!h2f_ARID_2),
	.datab(!h2f_AWID_2),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_107),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[107] .extended_lut = "off";
defparam \src_data[107] .lut_mask = 64'h0537053705370537;
defparam \src_data[107] .shared_arith = "off";

cyclonev_lcell_comb \src_data[108] (
	.dataa(!h2f_ARID_3),
	.datab(!h2f_AWID_3),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_108),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[108] .extended_lut = "off";
defparam \src_data[108] .lut_mask = 64'h0537053705370537;
defparam \src_data[108] .shared_arith = "off";

cyclonev_lcell_comb \src_data[109] (
	.dataa(!h2f_ARID_4),
	.datab(!h2f_AWID_4),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_109),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[109] .extended_lut = "off";
defparam \src_data[109] .lut_mask = 64'h0537053705370537;
defparam \src_data[109] .shared_arith = "off";

cyclonev_lcell_comb \src_data[110] (
	.dataa(!h2f_ARID_5),
	.datab(!h2f_AWID_5),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_110),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[110] .extended_lut = "off";
defparam \src_data[110] .lut_mask = 64'h0537053705370537;
defparam \src_data[110] .shared_arith = "off";

cyclonev_lcell_comb \src_data[111] (
	.dataa(!h2f_ARID_6),
	.datab(!h2f_AWID_6),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_111),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[111] .extended_lut = "off";
defparam \src_data[111] .lut_mask = 64'h0537053705370537;
defparam \src_data[111] .shared_arith = "off";

cyclonev_lcell_comb \src_data[112] (
	.dataa(!h2f_ARID_7),
	.datab(!h2f_AWID_7),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_112),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[112] .extended_lut = "off";
defparam \src_data[112] .lut_mask = 64'h0537053705370537;
defparam \src_data[112] .shared_arith = "off";

cyclonev_lcell_comb \src_data[113] (
	.dataa(!h2f_ARID_8),
	.datab(!h2f_AWID_8),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_113),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[113] .extended_lut = "off";
defparam \src_data[113] .lut_mask = 64'h0537053705370537;
defparam \src_data[113] .shared_arith = "off";

cyclonev_lcell_comb \src_data[114] (
	.dataa(!h2f_ARID_9),
	.datab(!h2f_AWID_9),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_114),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[114] .extended_lut = "off";
defparam \src_data[114] .lut_mask = 64'h0537053705370537;
defparam \src_data[114] .shared_arith = "off";

cyclonev_lcell_comb \src_data[115] (
	.dataa(!h2f_ARID_10),
	.datab(!h2f_AWID_10),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_115),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[115] .extended_lut = "off";
defparam \src_data[115] .lut_mask = 64'h0537053705370537;
defparam \src_data[115] .shared_arith = "off";

cyclonev_lcell_comb \src_data[116] (
	.dataa(!h2f_ARID_11),
	.datab(!h2f_AWID_11),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_116),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[116] .extended_lut = "off";
defparam \src_data[116] .lut_mask = 64'h0537053705370537;
defparam \src_data[116] .shared_arith = "off";

cyclonev_lcell_comb \src_data[86] (
	.dataa(!h2f_ARSIZE_0),
	.datab(!h2f_AWSIZE_0),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_86),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[86] .extended_lut = "off";
defparam \src_data[86] .lut_mask = 64'h0537053705370537;
defparam \src_data[86] .shared_arith = "off";

cyclonev_lcell_comb \src_data[80] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector5),
	.datad(!Selector12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_80),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[80] .extended_lut = "off";
defparam \src_data[80] .lut_mask = 64'h0357035703570357;
defparam \src_data[80] .shared_arith = "off";

cyclonev_lcell_comb \src_data[79] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector6),
	.datad(!Selector13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_79),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[79] .extended_lut = "off";
defparam \src_data[79] .lut_mask = 64'h0357035703570357;
defparam \src_data[79] .shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!\update_grant~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \update_grant~0 (
	.dataa(!nxt_in_ready1),
	.datab(!nxt_in_ready),
	.datac(!src_valid),
	.datad(!src_valid1),
	.datae(!src_payload_0),
	.dataf(!\packet_in_progress~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\update_grant~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \update_grant~0 .extended_lut = "off";
defparam \update_grant~0 .lut_mask = 64'hF000F77700000777;
defparam \update_grant~0 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_arbitrator_1 (
	nxt_in_ready,
	nxt_in_ready1,
	Equal16,
	reset,
	Equal14,
	src2_valid,
	src_payload_0,
	src2_valid1,
	src2_valid2,
	grant_1,
	packet_in_progress,
	grant_0,
	WideOr1,
	clk)/* synthesis synthesis_greybox=0 */;
input 	nxt_in_ready;
input 	nxt_in_ready1;
input 	Equal16;
input 	reset;
input 	Equal14;
input 	src2_valid;
input 	src_payload_0;
input 	src2_valid1;
input 	src2_valid2;
output 	grant_1;
input 	packet_in_progress;
output 	grant_0;
input 	WideOr1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg[0]~2_combout ;
wire \top_priority_reg[0]~q ;


cyclonev_lcell_comb \grant[1]~0 (
	.dataa(!\top_priority_reg[1]~q ),
	.datab(!\top_priority_reg[0]~q ),
	.datac(!src2_valid1),
	.datad(!src2_valid2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[1]~0 .extended_lut = "off";
defparam \grant[1]~0 .lut_mask = 64'h00D500D500D500D5;
defparam \grant[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \grant[0]~1 (
	.dataa(!\top_priority_reg[1]~q ),
	.datab(!\top_priority_reg[0]~q ),
	.datac(!src2_valid1),
	.datad(!src2_valid2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[0]~1 .extended_lut = "off";
defparam \grant[0]~1 .lut_mask = 64'h0D0C0D0C0D0C0D0C;
defparam \grant[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~0 (
	.dataa(!Equal16),
	.datab(!Equal14),
	.datac(!src2_valid),
	.datad(!src2_valid2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~0 .extended_lut = "off";
defparam \top_priority_reg[0]~0 .lut_mask = 64'hFE00FE00FE00FE00;
defparam \top_priority_reg[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~1 (
	.dataa(!nxt_in_ready1),
	.datab(!nxt_in_ready),
	.datac(!WideOr1),
	.datad(!src_payload_0),
	.datae(!packet_in_progress),
	.dataf(!\top_priority_reg[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~1 .extended_lut = "off";
defparam \top_priority_reg[0]~1 .lut_mask = 64'h0F7F007000000000;
defparam \top_priority_reg[0]~1 .shared_arith = "off";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~1_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

cyclonev_lcell_comb \top_priority_reg[0]~2 (
	.dataa(!grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~2 .extended_lut = "off";
defparam \top_priority_reg[0]~2 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \top_priority_reg[0]~2 .shared_arith = "off";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~1_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

endmodule

module spw_babasu_spw_babasu_mm_interconnect_0_cmd_mux_3 (
	h2f_ARVALID_0,
	h2f_ARSIZE_0,
	h2f_ARSIZE_1,
	h2f_ARSIZE_2,
	has_pending_responses,
	Equal3,
	saved_grant_1,
	altera_reset_synchronizer_int_chain_out,
	nxt_in_ready,
	last_channel_3,
	src_valid,
	src_payload,
	src_payload1,
	src_payload2,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARVALID_0;
input 	h2f_ARSIZE_0;
input 	h2f_ARSIZE_1;
input 	h2f_ARSIZE_2;
input 	has_pending_responses;
input 	Equal3;
output 	saved_grant_1;
input 	altera_reset_synchronizer_int_chain_out;
input 	nxt_in_ready;
input 	last_channel_3;
output 	src_valid;
output 	src_payload;
output 	src_payload1;
output 	src_payload2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \last_cycle~0_combout ;
wire \saved_grant[1]~0_combout ;


dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\saved_grant[1]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cyclonev_lcell_comb \src_valid~0 (
	.dataa(!saved_grant_1),
	.datab(!\last_cycle~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~0 .extended_lut = "off";
defparam \src_valid~0 .lut_mask = 64'h1111111111111111;
defparam \src_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!h2f_ARSIZE_0),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h1111111111111111;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!h2f_ARSIZE_2),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h1111111111111111;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!h2f_ARSIZE_1),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h1111111111111111;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!nxt_in_ready),
	.datab(!\packet_in_progress~q ),
	.datac(!src_valid),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'h3535353535353535;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \last_cycle~0 (
	.dataa(!h2f_ARVALID_0),
	.datab(!has_pending_responses),
	.datac(!Equal3),
	.datad(!last_channel_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_cycle~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_cycle~0 .extended_lut = "off";
defparam \last_cycle~0 .lut_mask = 64'h0405040504050405;
defparam \last_cycle~0 .shared_arith = "off";

cyclonev_lcell_comb \saved_grant[1]~0 (
	.dataa(!saved_grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(!\packet_in_progress~q ),
	.datae(!\last_cycle~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\saved_grant[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \saved_grant[1]~0 .extended_lut = "off";
defparam \saved_grant[1]~0 .lut_mask = 64'h0055FF550055FF55;
defparam \saved_grant[1]~0 .shared_arith = "off";

endmodule

module spw_babasu_spw_babasu_mm_interconnect_0_cmd_mux_4 (
	h2f_ARVALID_0,
	h2f_ARSIZE_0,
	h2f_ARSIZE_1,
	h2f_ARSIZE_2,
	has_pending_responses,
	saved_grant_1,
	altera_reset_synchronizer_int_chain_out,
	nxt_in_ready,
	Equal4,
	last_channel_4,
	src_valid,
	src_payload,
	src_payload1,
	src_payload2,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARVALID_0;
input 	h2f_ARSIZE_0;
input 	h2f_ARSIZE_1;
input 	h2f_ARSIZE_2;
input 	has_pending_responses;
output 	saved_grant_1;
input 	altera_reset_synchronizer_int_chain_out;
input 	nxt_in_ready;
input 	Equal4;
input 	last_channel_4;
output 	src_valid;
output 	src_payload;
output 	src_payload1;
output 	src_payload2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \saved_grant[1]~0_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \saved_grant[1]~1_combout ;


dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\saved_grant[1]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cyclonev_lcell_comb \src_valid~0 (
	.dataa(!Equal4),
	.datab(!saved_grant_1),
	.datac(!\saved_grant[1]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~0 .extended_lut = "off";
defparam \src_valid~0 .lut_mask = 64'h0101010101010101;
defparam \src_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!h2f_ARSIZE_0),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h1111111111111111;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!h2f_ARSIZE_2),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h1111111111111111;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!h2f_ARSIZE_1),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h1111111111111111;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \saved_grant[1]~0 (
	.dataa(!h2f_ARVALID_0),
	.datab(!has_pending_responses),
	.datac(!last_channel_4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\saved_grant[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \saved_grant[1]~0 .extended_lut = "off";
defparam \saved_grant[1]~0 .lut_mask = 64'h4545454545454545;
defparam \saved_grant[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!nxt_in_ready),
	.datab(!\packet_in_progress~q ),
	.datac(!src_valid),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'h3535353535353535;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \saved_grant[1]~1 (
	.dataa(!Equal4),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(!\saved_grant[1]~0_combout ),
	.datae(!\packet_in_progress~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\saved_grant[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \saved_grant[1]~1 .extended_lut = "off";
defparam \saved_grant[1]~1 .lut_mask = 64'h0055333300553333;
defparam \saved_grant[1]~1 .shared_arith = "off";

endmodule

module spw_babasu_spw_babasu_mm_interconnect_0_cmd_mux_5 (
	h2f_ARVALID_0,
	h2f_WLAST_0,
	h2f_ARADDR_4,
	h2f_ARADDR_5,
	h2f_ARADDR_6,
	h2f_ARADDR_7,
	h2f_ARADDR_8,
	h2f_ARID_0,
	h2f_ARID_1,
	h2f_ARID_2,
	h2f_ARID_3,
	h2f_ARID_4,
	h2f_ARID_5,
	h2f_ARID_6,
	h2f_ARID_7,
	h2f_ARID_8,
	h2f_ARID_9,
	h2f_ARID_10,
	h2f_ARID_11,
	h2f_ARSIZE_0,
	h2f_ARSIZE_1,
	h2f_ARSIZE_2,
	h2f_AWID_0,
	h2f_AWID_1,
	h2f_AWID_2,
	h2f_AWID_3,
	h2f_AWID_4,
	h2f_AWID_5,
	h2f_AWID_6,
	h2f_AWID_7,
	h2f_AWID_8,
	h2f_AWID_9,
	h2f_AWID_10,
	h2f_AWID_11,
	h2f_AWSIZE_0,
	h2f_AWSIZE_1,
	h2f_AWSIZE_2,
	h2f_WDATA_0,
	h2f_WDATA_1,
	h2f_WDATA_2,
	h2f_WDATA_3,
	h2f_WDATA_4,
	h2f_WDATA_5,
	h2f_WDATA_6,
	h2f_WDATA_7,
	h2f_WDATA_8,
	h2f_WSTRB_0,
	h2f_WSTRB_1,
	h2f_WSTRB_2,
	h2f_WSTRB_3,
	nxt_in_ready,
	nxt_in_ready1,
	saved_grant_1,
	write_addr_data_both_valid,
	out_data_5,
	Equal5,
	Equal15,
	saved_grant_0,
	altera_reset_synchronizer_int_chain_out,
	Equal51,
	src5_valid,
	src5_valid1,
	cmd_src_valid_5,
	src_valid,
	src_data_87,
	src_data_88,
	src_valid1,
	src_data_35,
	src_data_34,
	src_data_33,
	src_data_32,
	src_payload_0,
	src5_valid2,
	Selector3,
	Selector10,
	Selector4,
	Selector11,
	src_payload,
	src_data_82,
	src_data_81,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_data_105,
	src_data_106,
	src_data_107,
	src_data_108,
	src_data_109,
	src_data_110,
	src_data_111,
	src_data_112,
	src_data_113,
	src_data_114,
	src_data_115,
	src_data_116,
	src_data_86,
	Selector5,
	Selector12,
	src_data_80,
	Selector6,
	Selector13,
	src_data_79,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARVALID_0;
input 	h2f_WLAST_0;
input 	h2f_ARADDR_4;
input 	h2f_ARADDR_5;
input 	h2f_ARADDR_6;
input 	h2f_ARADDR_7;
input 	h2f_ARADDR_8;
input 	h2f_ARID_0;
input 	h2f_ARID_1;
input 	h2f_ARID_2;
input 	h2f_ARID_3;
input 	h2f_ARID_4;
input 	h2f_ARID_5;
input 	h2f_ARID_6;
input 	h2f_ARID_7;
input 	h2f_ARID_8;
input 	h2f_ARID_9;
input 	h2f_ARID_10;
input 	h2f_ARID_11;
input 	h2f_ARSIZE_0;
input 	h2f_ARSIZE_1;
input 	h2f_ARSIZE_2;
input 	h2f_AWID_0;
input 	h2f_AWID_1;
input 	h2f_AWID_2;
input 	h2f_AWID_3;
input 	h2f_AWID_4;
input 	h2f_AWID_5;
input 	h2f_AWID_6;
input 	h2f_AWID_7;
input 	h2f_AWID_8;
input 	h2f_AWID_9;
input 	h2f_AWID_10;
input 	h2f_AWID_11;
input 	h2f_AWSIZE_0;
input 	h2f_AWSIZE_1;
input 	h2f_AWSIZE_2;
input 	h2f_WDATA_0;
input 	h2f_WDATA_1;
input 	h2f_WDATA_2;
input 	h2f_WDATA_3;
input 	h2f_WDATA_4;
input 	h2f_WDATA_5;
input 	h2f_WDATA_6;
input 	h2f_WDATA_7;
input 	h2f_WDATA_8;
input 	h2f_WSTRB_0;
input 	h2f_WSTRB_1;
input 	h2f_WSTRB_2;
input 	h2f_WSTRB_3;
input 	nxt_in_ready;
input 	nxt_in_ready1;
output 	saved_grant_1;
input 	write_addr_data_both_valid;
input 	out_data_5;
input 	Equal5;
input 	Equal15;
output 	saved_grant_0;
input 	altera_reset_synchronizer_int_chain_out;
input 	Equal51;
input 	src5_valid;
input 	src5_valid1;
input 	cmd_src_valid_5;
output 	src_valid;
output 	src_data_87;
output 	src_data_88;
output 	src_valid1;
output 	src_data_35;
output 	src_data_34;
output 	src_data_33;
output 	src_data_32;
output 	src_payload_0;
input 	src5_valid2;
input 	Selector3;
input 	Selector10;
input 	Selector4;
input 	Selector11;
output 	src_payload;
output 	src_data_82;
output 	src_data_81;
output 	src_payload1;
output 	src_payload2;
output 	src_payload3;
output 	src_payload4;
output 	src_payload5;
output 	src_payload6;
output 	src_payload7;
output 	src_payload8;
output 	src_data_105;
output 	src_data_106;
output 	src_data_107;
output 	src_data_108;
output 	src_data_109;
output 	src_data_110;
output 	src_data_111;
output 	src_data_112;
output 	src_data_113;
output 	src_data_114;
output 	src_data_115;
output 	src_data_116;
output 	src_data_86;
input 	Selector5;
input 	Selector12;
output 	src_data_80;
input 	Selector6;
input 	Selector13;
output 	src_data_79;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \src_valid~3_combout ;
wire \arb|grant[1]~0_combout ;
wire \arb|grant[0]~1_combout ;
wire \WideOr1~combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~0_combout ;
wire \src_valid~0_combout ;


spw_babasu_altera_merlin_arbitrator_4 arb(
	.nxt_in_ready(nxt_in_ready),
	.nxt_in_ready1(nxt_in_ready1),
	.Equal5(Equal5),
	.reset(altera_reset_synchronizer_int_chain_out),
	.Equal51(Equal51),
	.src5_valid(src5_valid1),
	.src_payload_0(src_payload_0),
	.src5_valid1(src5_valid2),
	.src_valid(\src_valid~3_combout ),
	.grant_1(\arb|grant[1]~0_combout ),
	.packet_in_progress(\packet_in_progress~q ),
	.grant_0(\arb|grant[0]~1_combout ),
	.WideOr1(\WideOr1~combout ),
	.clk(clk_clk));

cyclonev_lcell_comb \src_valid~3 (
	.dataa(!cmd_src_valid_5),
	.datab(!\src_valid~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_valid~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~3 .extended_lut = "off";
defparam \src_valid~3 .lut_mask = 64'h2222222222222222;
defparam \src_valid~3 .shared_arith = "off";

cyclonev_lcell_comb WideOr1(
	.dataa(!Equal51),
	.datab(!Equal5),
	.datac(!saved_grant_0),
	.datad(!src5_valid1),
	.datae(!src_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr1.extended_lut = "off";
defparam WideOr1.lut_mask = 64'hFFFE0000FFFE0000;
defparam WideOr1.shared_arith = "off";

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

cyclonev_lcell_comb \src_valid~1 (
	.dataa(!saved_grant_1),
	.datab(!cmd_src_valid_5),
	.datac(!\src_valid~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~1 .extended_lut = "off";
defparam \src_valid~1 .lut_mask = 64'h0404040404040404;
defparam \src_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \src_data[87] (
	.dataa(!h2f_ARSIZE_1),
	.datab(!h2f_AWSIZE_1),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_87),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[87] .extended_lut = "off";
defparam \src_data[87] .lut_mask = 64'h0537053705370537;
defparam \src_data[87] .shared_arith = "off";

cyclonev_lcell_comb \src_data[88] (
	.dataa(!h2f_ARSIZE_2),
	.datab(!h2f_AWSIZE_2),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_88),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[88] .extended_lut = "off";
defparam \src_data[88] .lut_mask = 64'h0537053705370537;
defparam \src_data[88] .shared_arith = "off";

cyclonev_lcell_comb \src_valid~2 (
	.dataa(!out_data_5),
	.datab(!Equal15),
	.datac(!Equal5),
	.datad(!saved_grant_0),
	.datae(!write_addr_data_both_valid),
	.dataf(!src5_valid),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~2 .extended_lut = "off";
defparam \src_valid~2 .lut_mask = 64'h0000000200000000;
defparam \src_valid~2 .shared_arith = "off";

cyclonev_lcell_comb \src_data[35] (
	.dataa(!h2f_WSTRB_3),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_35),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[35] .extended_lut = "off";
defparam \src_data[35] .lut_mask = 64'h3737373737373737;
defparam \src_data[35] .shared_arith = "off";

cyclonev_lcell_comb \src_data[34] (
	.dataa(!h2f_WSTRB_2),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_34),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[34] .extended_lut = "off";
defparam \src_data[34] .lut_mask = 64'h3737373737373737;
defparam \src_data[34] .shared_arith = "off";

cyclonev_lcell_comb \src_data[33] (
	.dataa(!h2f_WSTRB_1),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_33),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[33] .extended_lut = "off";
defparam \src_data[33] .lut_mask = 64'h3737373737373737;
defparam \src_data[33] .shared_arith = "off";

cyclonev_lcell_comb \src_data[32] (
	.dataa(!h2f_WSTRB_0),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_32),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[32] .extended_lut = "off";
defparam \src_data[32] .lut_mask = 64'h3737373737373737;
defparam \src_data[32] .shared_arith = "off";

cyclonev_lcell_comb \src_payload[0] (
	.dataa(!h2f_WLAST_0),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload[0] .extended_lut = "off";
defparam \src_payload[0] .lut_mask = 64'h3737373737373737;
defparam \src_payload[0] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!h2f_WDATA_0),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h1111111111111111;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[82] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector3),
	.datad(!Selector10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_82),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[82] .extended_lut = "off";
defparam \src_data[82] .lut_mask = 64'h0357035703570357;
defparam \src_data[82] .shared_arith = "off";

cyclonev_lcell_comb \src_data[81] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector4),
	.datad(!Selector11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_81),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[81] .extended_lut = "off";
defparam \src_data[81] .lut_mask = 64'h0357035703570357;
defparam \src_data[81] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!h2f_WDATA_1),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h1111111111111111;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!h2f_WDATA_2),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h1111111111111111;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~3 (
	.dataa(!h2f_WDATA_3),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~3 .extended_lut = "off";
defparam \src_payload~3 .lut_mask = 64'h1111111111111111;
defparam \src_payload~3 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~4 (
	.dataa(!h2f_WDATA_4),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~4 .extended_lut = "off";
defparam \src_payload~4 .lut_mask = 64'h1111111111111111;
defparam \src_payload~4 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~5 (
	.dataa(!h2f_WDATA_5),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~5 .extended_lut = "off";
defparam \src_payload~5 .lut_mask = 64'h1111111111111111;
defparam \src_payload~5 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~6 (
	.dataa(!h2f_WDATA_6),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~6 .extended_lut = "off";
defparam \src_payload~6 .lut_mask = 64'h1111111111111111;
defparam \src_payload~6 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~7 (
	.dataa(!h2f_WDATA_7),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~7 .extended_lut = "off";
defparam \src_payload~7 .lut_mask = 64'h1111111111111111;
defparam \src_payload~7 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~8 (
	.dataa(!h2f_WDATA_8),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~8 .extended_lut = "off";
defparam \src_payload~8 .lut_mask = 64'h1111111111111111;
defparam \src_payload~8 .shared_arith = "off";

cyclonev_lcell_comb \src_data[105] (
	.dataa(!h2f_ARID_0),
	.datab(!h2f_AWID_0),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_105),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[105] .extended_lut = "off";
defparam \src_data[105] .lut_mask = 64'h0537053705370537;
defparam \src_data[105] .shared_arith = "off";

cyclonev_lcell_comb \src_data[106] (
	.dataa(!h2f_ARID_1),
	.datab(!h2f_AWID_1),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_106),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[106] .extended_lut = "off";
defparam \src_data[106] .lut_mask = 64'h0537053705370537;
defparam \src_data[106] .shared_arith = "off";

cyclonev_lcell_comb \src_data[107] (
	.dataa(!h2f_ARID_2),
	.datab(!h2f_AWID_2),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_107),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[107] .extended_lut = "off";
defparam \src_data[107] .lut_mask = 64'h0537053705370537;
defparam \src_data[107] .shared_arith = "off";

cyclonev_lcell_comb \src_data[108] (
	.dataa(!h2f_ARID_3),
	.datab(!h2f_AWID_3),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_108),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[108] .extended_lut = "off";
defparam \src_data[108] .lut_mask = 64'h0537053705370537;
defparam \src_data[108] .shared_arith = "off";

cyclonev_lcell_comb \src_data[109] (
	.dataa(!h2f_ARID_4),
	.datab(!h2f_AWID_4),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_109),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[109] .extended_lut = "off";
defparam \src_data[109] .lut_mask = 64'h0537053705370537;
defparam \src_data[109] .shared_arith = "off";

cyclonev_lcell_comb \src_data[110] (
	.dataa(!h2f_ARID_5),
	.datab(!h2f_AWID_5),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_110),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[110] .extended_lut = "off";
defparam \src_data[110] .lut_mask = 64'h0537053705370537;
defparam \src_data[110] .shared_arith = "off";

cyclonev_lcell_comb \src_data[111] (
	.dataa(!h2f_ARID_6),
	.datab(!h2f_AWID_6),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_111),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[111] .extended_lut = "off";
defparam \src_data[111] .lut_mask = 64'h0537053705370537;
defparam \src_data[111] .shared_arith = "off";

cyclonev_lcell_comb \src_data[112] (
	.dataa(!h2f_ARID_7),
	.datab(!h2f_AWID_7),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_112),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[112] .extended_lut = "off";
defparam \src_data[112] .lut_mask = 64'h0537053705370537;
defparam \src_data[112] .shared_arith = "off";

cyclonev_lcell_comb \src_data[113] (
	.dataa(!h2f_ARID_8),
	.datab(!h2f_AWID_8),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_113),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[113] .extended_lut = "off";
defparam \src_data[113] .lut_mask = 64'h0537053705370537;
defparam \src_data[113] .shared_arith = "off";

cyclonev_lcell_comb \src_data[114] (
	.dataa(!h2f_ARID_9),
	.datab(!h2f_AWID_9),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_114),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[114] .extended_lut = "off";
defparam \src_data[114] .lut_mask = 64'h0537053705370537;
defparam \src_data[114] .shared_arith = "off";

cyclonev_lcell_comb \src_data[115] (
	.dataa(!h2f_ARID_10),
	.datab(!h2f_AWID_10),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_115),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[115] .extended_lut = "off";
defparam \src_data[115] .lut_mask = 64'h0537053705370537;
defparam \src_data[115] .shared_arith = "off";

cyclonev_lcell_comb \src_data[116] (
	.dataa(!h2f_ARID_11),
	.datab(!h2f_AWID_11),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_116),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[116] .extended_lut = "off";
defparam \src_data[116] .lut_mask = 64'h0537053705370537;
defparam \src_data[116] .shared_arith = "off";

cyclonev_lcell_comb \src_data[86] (
	.dataa(!h2f_ARSIZE_0),
	.datab(!h2f_AWSIZE_0),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_86),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[86] .extended_lut = "off";
defparam \src_data[86] .lut_mask = 64'h0537053705370537;
defparam \src_data[86] .shared_arith = "off";

cyclonev_lcell_comb \src_data[80] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector5),
	.datad(!Selector12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_80),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[80] .extended_lut = "off";
defparam \src_data[80] .lut_mask = 64'h0357035703570357;
defparam \src_data[80] .shared_arith = "off";

cyclonev_lcell_comb \src_data[79] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector6),
	.datad(!Selector13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_79),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[79] .extended_lut = "off";
defparam \src_data[79] .lut_mask = 64'h0357035703570357;
defparam \src_data[79] .shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!\update_grant~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \update_grant~0 (
	.dataa(!nxt_in_ready1),
	.datab(!nxt_in_ready),
	.datac(!src_valid),
	.datad(!src_valid1),
	.datae(!src_payload_0),
	.dataf(!\packet_in_progress~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\update_grant~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \update_grant~0 .extended_lut = "off";
defparam \update_grant~0 .lut_mask = 64'hF000F77700000777;
defparam \update_grant~0 .shared_arith = "off";

cyclonev_lcell_comb \src_valid~0 (
	.dataa(!h2f_ARVALID_0),
	.datab(!h2f_ARADDR_4),
	.datac(!h2f_ARADDR_5),
	.datad(!h2f_ARADDR_6),
	.datae(!h2f_ARADDR_7),
	.dataf(!h2f_ARADDR_8),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~0 .extended_lut = "off";
defparam \src_valid~0 .lut_mask = 64'h0010000000000000;
defparam \src_valid~0 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_arbitrator_4 (
	nxt_in_ready,
	nxt_in_ready1,
	Equal5,
	reset,
	Equal51,
	src5_valid,
	src_payload_0,
	src5_valid1,
	src_valid,
	grant_1,
	packet_in_progress,
	grant_0,
	WideOr1,
	clk)/* synthesis synthesis_greybox=0 */;
input 	nxt_in_ready;
input 	nxt_in_ready1;
input 	Equal5;
input 	reset;
input 	Equal51;
input 	src5_valid;
input 	src_payload_0;
input 	src5_valid1;
input 	src_valid;
output 	grant_1;
input 	packet_in_progress;
output 	grant_0;
input 	WideOr1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg[0]~2_combout ;
wire \top_priority_reg[0]~q ;


cyclonev_lcell_comb \grant[1]~0 (
	.dataa(!\top_priority_reg[1]~q ),
	.datab(!\top_priority_reg[0]~q ),
	.datac(!src5_valid1),
	.datad(!src_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[1]~0 .extended_lut = "off";
defparam \grant[1]~0 .lut_mask = 64'h00D500D500D500D5;
defparam \grant[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \grant[0]~1 (
	.dataa(!\top_priority_reg[1]~q ),
	.datab(!\top_priority_reg[0]~q ),
	.datac(!src5_valid1),
	.datad(!src_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[0]~1 .extended_lut = "off";
defparam \grant[0]~1 .lut_mask = 64'h0D0C0D0C0D0C0D0C;
defparam \grant[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~0 (
	.dataa(!Equal51),
	.datab(!Equal5),
	.datac(!src5_valid),
	.datad(!src_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~0 .extended_lut = "off";
defparam \top_priority_reg[0]~0 .lut_mask = 64'hFE00FE00FE00FE00;
defparam \top_priority_reg[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~1 (
	.dataa(!nxt_in_ready1),
	.datab(!nxt_in_ready),
	.datac(!WideOr1),
	.datad(!src_payload_0),
	.datae(!packet_in_progress),
	.dataf(!\top_priority_reg[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~1 .extended_lut = "off";
defparam \top_priority_reg[0]~1 .lut_mask = 64'h0F7F007000000000;
defparam \top_priority_reg[0]~1 .shared_arith = "off";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~1_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

cyclonev_lcell_comb \top_priority_reg[0]~2 (
	.dataa(!grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~2 .extended_lut = "off";
defparam \top_priority_reg[0]~2 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \top_priority_reg[0]~2 .shared_arith = "off";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~1_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

endmodule

module spw_babasu_spw_babasu_mm_interconnect_0_cmd_mux_6 (
	h2f_WLAST_0,
	h2f_ARID_0,
	h2f_ARID_1,
	h2f_ARID_2,
	h2f_ARID_3,
	h2f_ARID_4,
	h2f_ARID_5,
	h2f_ARID_6,
	h2f_ARID_7,
	h2f_ARID_8,
	h2f_ARID_9,
	h2f_ARID_10,
	h2f_ARID_11,
	h2f_ARSIZE_0,
	h2f_ARSIZE_1,
	h2f_ARSIZE_2,
	h2f_AWID_0,
	h2f_AWID_1,
	h2f_AWID_2,
	h2f_AWID_3,
	h2f_AWID_4,
	h2f_AWID_5,
	h2f_AWID_6,
	h2f_AWID_7,
	h2f_AWID_8,
	h2f_AWID_9,
	h2f_AWID_10,
	h2f_AWID_11,
	h2f_AWSIZE_0,
	h2f_AWSIZE_1,
	h2f_AWSIZE_2,
	h2f_WDATA_0,
	h2f_WSTRB_0,
	h2f_WSTRB_1,
	h2f_WSTRB_2,
	h2f_WSTRB_3,
	nxt_in_ready,
	Equal6,
	nxt_in_ready1,
	saved_grant_1,
	write_addr_data_both_valid,
	out_data_4,
	Equal5,
	Equal14,
	saved_grant_0,
	altera_reset_synchronizer_int_chain_out,
	Equal141,
	src6_valid,
	src6_valid1,
	src6_valid2,
	src_valid,
	src_data_87,
	src_data_88,
	src_valid1,
	src_data_35,
	src_data_34,
	src_data_33,
	src_data_32,
	src_payload_0,
	src6_valid3,
	src6_valid4,
	Selector3,
	Selector10,
	Selector4,
	Selector11,
	src_payload,
	src_data_82,
	src_data_81,
	src_data_105,
	src_data_106,
	src_data_107,
	src_data_108,
	src_data_109,
	src_data_110,
	src_data_111,
	src_data_112,
	src_data_113,
	src_data_114,
	src_data_115,
	src_data_116,
	src_data_86,
	Selector5,
	Selector12,
	src_data_80,
	Selector6,
	Selector13,
	src_data_79,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_WLAST_0;
input 	h2f_ARID_0;
input 	h2f_ARID_1;
input 	h2f_ARID_2;
input 	h2f_ARID_3;
input 	h2f_ARID_4;
input 	h2f_ARID_5;
input 	h2f_ARID_6;
input 	h2f_ARID_7;
input 	h2f_ARID_8;
input 	h2f_ARID_9;
input 	h2f_ARID_10;
input 	h2f_ARID_11;
input 	h2f_ARSIZE_0;
input 	h2f_ARSIZE_1;
input 	h2f_ARSIZE_2;
input 	h2f_AWID_0;
input 	h2f_AWID_1;
input 	h2f_AWID_2;
input 	h2f_AWID_3;
input 	h2f_AWID_4;
input 	h2f_AWID_5;
input 	h2f_AWID_6;
input 	h2f_AWID_7;
input 	h2f_AWID_8;
input 	h2f_AWID_9;
input 	h2f_AWID_10;
input 	h2f_AWID_11;
input 	h2f_AWSIZE_0;
input 	h2f_AWSIZE_1;
input 	h2f_AWSIZE_2;
input 	h2f_WDATA_0;
input 	h2f_WSTRB_0;
input 	h2f_WSTRB_1;
input 	h2f_WSTRB_2;
input 	h2f_WSTRB_3;
input 	nxt_in_ready;
input 	Equal6;
input 	nxt_in_ready1;
output 	saved_grant_1;
input 	write_addr_data_both_valid;
input 	out_data_4;
input 	Equal5;
input 	Equal14;
output 	saved_grant_0;
input 	altera_reset_synchronizer_int_chain_out;
input 	Equal141;
input 	src6_valid;
input 	src6_valid1;
input 	src6_valid2;
output 	src_valid;
output 	src_data_87;
output 	src_data_88;
output 	src_valid1;
output 	src_data_35;
output 	src_data_34;
output 	src_data_33;
output 	src_data_32;
output 	src_payload_0;
input 	src6_valid3;
input 	src6_valid4;
input 	Selector3;
input 	Selector10;
input 	Selector4;
input 	Selector11;
output 	src_payload;
output 	src_data_82;
output 	src_data_81;
output 	src_data_105;
output 	src_data_106;
output 	src_data_107;
output 	src_data_108;
output 	src_data_109;
output 	src_data_110;
output 	src_data_111;
output 	src_data_112;
output 	src_data_113;
output 	src_data_114;
output 	src_data_115;
output 	src_data_116;
output 	src_data_86;
input 	Selector5;
input 	Selector12;
output 	src_data_80;
input 	Selector6;
input 	Selector13;
output 	src_data_79;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[1]~0_combout ;
wire \arb|grant[0]~1_combout ;
wire \WideOr1~combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~0_combout ;


spw_babasu_altera_merlin_arbitrator_5 arb(
	.nxt_in_ready(nxt_in_ready),
	.nxt_in_ready1(nxt_in_ready1),
	.Equal5(Equal5),
	.reset(altera_reset_synchronizer_int_chain_out),
	.Equal14(Equal141),
	.src6_valid(src6_valid1),
	.src_payload_0(src_payload_0),
	.src6_valid1(src6_valid3),
	.src6_valid2(src6_valid4),
	.grant_1(\arb|grant[1]~0_combout ),
	.packet_in_progress(\packet_in_progress~q ),
	.grant_0(\arb|grant[0]~1_combout ),
	.WideOr1(\WideOr1~combout ),
	.clk(clk_clk));

cyclonev_lcell_comb WideOr1(
	.dataa(!Equal5),
	.datab(!Equal141),
	.datac(!saved_grant_0),
	.datad(!src6_valid1),
	.datae(!src_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr1.extended_lut = "off";
defparam WideOr1.lut_mask = 64'hFFFE0000FFFE0000;
defparam WideOr1.shared_arith = "off";

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

cyclonev_lcell_comb \src_valid~0 (
	.dataa(!Equal6),
	.datab(!saved_grant_1),
	.datac(!src6_valid2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~0 .extended_lut = "off";
defparam \src_valid~0 .lut_mask = 64'h0101010101010101;
defparam \src_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[87] (
	.dataa(!h2f_ARSIZE_1),
	.datab(!h2f_AWSIZE_1),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_87),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[87] .extended_lut = "off";
defparam \src_data[87] .lut_mask = 64'h0537053705370537;
defparam \src_data[87] .shared_arith = "off";

cyclonev_lcell_comb \src_data[88] (
	.dataa(!h2f_ARSIZE_2),
	.datab(!h2f_AWSIZE_2),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_88),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[88] .extended_lut = "off";
defparam \src_data[88] .lut_mask = 64'h0537053705370537;
defparam \src_data[88] .shared_arith = "off";

cyclonev_lcell_comb \src_valid~1 (
	.dataa(!out_data_4),
	.datab(!Equal5),
	.datac(!Equal14),
	.datad(!saved_grant_0),
	.datae(!write_addr_data_both_valid),
	.dataf(!src6_valid),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~1 .extended_lut = "off";
defparam \src_valid~1 .lut_mask = 64'h0000000200000000;
defparam \src_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \src_data[35] (
	.dataa(!h2f_WSTRB_3),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_35),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[35] .extended_lut = "off";
defparam \src_data[35] .lut_mask = 64'h3737373737373737;
defparam \src_data[35] .shared_arith = "off";

cyclonev_lcell_comb \src_data[34] (
	.dataa(!h2f_WSTRB_2),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_34),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[34] .extended_lut = "off";
defparam \src_data[34] .lut_mask = 64'h3737373737373737;
defparam \src_data[34] .shared_arith = "off";

cyclonev_lcell_comb \src_data[33] (
	.dataa(!h2f_WSTRB_1),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_33),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[33] .extended_lut = "off";
defparam \src_data[33] .lut_mask = 64'h3737373737373737;
defparam \src_data[33] .shared_arith = "off";

cyclonev_lcell_comb \src_data[32] (
	.dataa(!h2f_WSTRB_0),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_32),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[32] .extended_lut = "off";
defparam \src_data[32] .lut_mask = 64'h3737373737373737;
defparam \src_data[32] .shared_arith = "off";

cyclonev_lcell_comb \src_payload[0] (
	.dataa(!h2f_WLAST_0),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload[0] .extended_lut = "off";
defparam \src_payload[0] .lut_mask = 64'h3737373737373737;
defparam \src_payload[0] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!h2f_WDATA_0),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h1111111111111111;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[82] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector3),
	.datad(!Selector10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_82),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[82] .extended_lut = "off";
defparam \src_data[82] .lut_mask = 64'h0357035703570357;
defparam \src_data[82] .shared_arith = "off";

cyclonev_lcell_comb \src_data[81] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector4),
	.datad(!Selector11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_81),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[81] .extended_lut = "off";
defparam \src_data[81] .lut_mask = 64'h0357035703570357;
defparam \src_data[81] .shared_arith = "off";

cyclonev_lcell_comb \src_data[105] (
	.dataa(!h2f_ARID_0),
	.datab(!h2f_AWID_0),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_105),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[105] .extended_lut = "off";
defparam \src_data[105] .lut_mask = 64'h0537053705370537;
defparam \src_data[105] .shared_arith = "off";

cyclonev_lcell_comb \src_data[106] (
	.dataa(!h2f_ARID_1),
	.datab(!h2f_AWID_1),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_106),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[106] .extended_lut = "off";
defparam \src_data[106] .lut_mask = 64'h0537053705370537;
defparam \src_data[106] .shared_arith = "off";

cyclonev_lcell_comb \src_data[107] (
	.dataa(!h2f_ARID_2),
	.datab(!h2f_AWID_2),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_107),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[107] .extended_lut = "off";
defparam \src_data[107] .lut_mask = 64'h0537053705370537;
defparam \src_data[107] .shared_arith = "off";

cyclonev_lcell_comb \src_data[108] (
	.dataa(!h2f_ARID_3),
	.datab(!h2f_AWID_3),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_108),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[108] .extended_lut = "off";
defparam \src_data[108] .lut_mask = 64'h0537053705370537;
defparam \src_data[108] .shared_arith = "off";

cyclonev_lcell_comb \src_data[109] (
	.dataa(!h2f_ARID_4),
	.datab(!h2f_AWID_4),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_109),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[109] .extended_lut = "off";
defparam \src_data[109] .lut_mask = 64'h0537053705370537;
defparam \src_data[109] .shared_arith = "off";

cyclonev_lcell_comb \src_data[110] (
	.dataa(!h2f_ARID_5),
	.datab(!h2f_AWID_5),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_110),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[110] .extended_lut = "off";
defparam \src_data[110] .lut_mask = 64'h0537053705370537;
defparam \src_data[110] .shared_arith = "off";

cyclonev_lcell_comb \src_data[111] (
	.dataa(!h2f_ARID_6),
	.datab(!h2f_AWID_6),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_111),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[111] .extended_lut = "off";
defparam \src_data[111] .lut_mask = 64'h0537053705370537;
defparam \src_data[111] .shared_arith = "off";

cyclonev_lcell_comb \src_data[112] (
	.dataa(!h2f_ARID_7),
	.datab(!h2f_AWID_7),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_112),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[112] .extended_lut = "off";
defparam \src_data[112] .lut_mask = 64'h0537053705370537;
defparam \src_data[112] .shared_arith = "off";

cyclonev_lcell_comb \src_data[113] (
	.dataa(!h2f_ARID_8),
	.datab(!h2f_AWID_8),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_113),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[113] .extended_lut = "off";
defparam \src_data[113] .lut_mask = 64'h0537053705370537;
defparam \src_data[113] .shared_arith = "off";

cyclonev_lcell_comb \src_data[114] (
	.dataa(!h2f_ARID_9),
	.datab(!h2f_AWID_9),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_114),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[114] .extended_lut = "off";
defparam \src_data[114] .lut_mask = 64'h0537053705370537;
defparam \src_data[114] .shared_arith = "off";

cyclonev_lcell_comb \src_data[115] (
	.dataa(!h2f_ARID_10),
	.datab(!h2f_AWID_10),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_115),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[115] .extended_lut = "off";
defparam \src_data[115] .lut_mask = 64'h0537053705370537;
defparam \src_data[115] .shared_arith = "off";

cyclonev_lcell_comb \src_data[116] (
	.dataa(!h2f_ARID_11),
	.datab(!h2f_AWID_11),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_116),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[116] .extended_lut = "off";
defparam \src_data[116] .lut_mask = 64'h0537053705370537;
defparam \src_data[116] .shared_arith = "off";

cyclonev_lcell_comb \src_data[86] (
	.dataa(!h2f_ARSIZE_0),
	.datab(!h2f_AWSIZE_0),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_86),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[86] .extended_lut = "off";
defparam \src_data[86] .lut_mask = 64'h0537053705370537;
defparam \src_data[86] .shared_arith = "off";

cyclonev_lcell_comb \src_data[80] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector5),
	.datad(!Selector12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_80),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[80] .extended_lut = "off";
defparam \src_data[80] .lut_mask = 64'h0357035703570357;
defparam \src_data[80] .shared_arith = "off";

cyclonev_lcell_comb \src_data[79] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector6),
	.datad(!Selector13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_79),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[79] .extended_lut = "off";
defparam \src_data[79] .lut_mask = 64'h0357035703570357;
defparam \src_data[79] .shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!\update_grant~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \update_grant~0 (
	.dataa(!nxt_in_ready1),
	.datab(!nxt_in_ready),
	.datac(!src_valid),
	.datad(!src_valid1),
	.datae(!src_payload_0),
	.dataf(!\packet_in_progress~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\update_grant~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \update_grant~0 .extended_lut = "off";
defparam \update_grant~0 .lut_mask = 64'hF000F77700000777;
defparam \update_grant~0 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_arbitrator_5 (
	nxt_in_ready,
	nxt_in_ready1,
	Equal5,
	reset,
	Equal14,
	src6_valid,
	src_payload_0,
	src6_valid1,
	src6_valid2,
	grant_1,
	packet_in_progress,
	grant_0,
	WideOr1,
	clk)/* synthesis synthesis_greybox=0 */;
input 	nxt_in_ready;
input 	nxt_in_ready1;
input 	Equal5;
input 	reset;
input 	Equal14;
input 	src6_valid;
input 	src_payload_0;
input 	src6_valid1;
input 	src6_valid2;
output 	grant_1;
input 	packet_in_progress;
output 	grant_0;
input 	WideOr1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg[0]~2_combout ;
wire \top_priority_reg[0]~q ;


cyclonev_lcell_comb \grant[1]~0 (
	.dataa(!\top_priority_reg[1]~q ),
	.datab(!\top_priority_reg[0]~q ),
	.datac(!src6_valid1),
	.datad(!src6_valid2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[1]~0 .extended_lut = "off";
defparam \grant[1]~0 .lut_mask = 64'h00D500D500D500D5;
defparam \grant[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \grant[0]~1 (
	.dataa(!\top_priority_reg[1]~q ),
	.datab(!\top_priority_reg[0]~q ),
	.datac(!src6_valid1),
	.datad(!src6_valid2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[0]~1 .extended_lut = "off";
defparam \grant[0]~1 .lut_mask = 64'h0D0C0D0C0D0C0D0C;
defparam \grant[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~0 (
	.dataa(!Equal5),
	.datab(!Equal14),
	.datac(!src6_valid),
	.datad(!src6_valid2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~0 .extended_lut = "off";
defparam \top_priority_reg[0]~0 .lut_mask = 64'hFE00FE00FE00FE00;
defparam \top_priority_reg[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~1 (
	.dataa(!nxt_in_ready1),
	.datab(!nxt_in_ready),
	.datac(!WideOr1),
	.datad(!src_payload_0),
	.datae(!packet_in_progress),
	.dataf(!\top_priority_reg[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~1 .extended_lut = "off";
defparam \top_priority_reg[0]~1 .lut_mask = 64'h0F7F007000000000;
defparam \top_priority_reg[0]~1 .shared_arith = "off";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~1_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

cyclonev_lcell_comb \top_priority_reg[0]~2 (
	.dataa(!grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~2 .extended_lut = "off";
defparam \top_priority_reg[0]~2 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \top_priority_reg[0]~2 .shared_arith = "off";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~1_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

endmodule

module spw_babasu_spw_babasu_mm_interconnect_0_cmd_mux_7 (
	h2f_ARVALID_0,
	h2f_ARSIZE_0,
	h2f_ARSIZE_1,
	h2f_ARSIZE_2,
	has_pending_responses,
	saved_grant_1,
	altera_reset_synchronizer_int_chain_out,
	nxt_in_ready,
	Equal7,
	last_channel_7,
	src_valid,
	src_payload,
	src_payload1,
	src_payload2,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARVALID_0;
input 	h2f_ARSIZE_0;
input 	h2f_ARSIZE_1;
input 	h2f_ARSIZE_2;
input 	has_pending_responses;
output 	saved_grant_1;
input 	altera_reset_synchronizer_int_chain_out;
input 	nxt_in_ready;
input 	Equal7;
input 	last_channel_7;
output 	src_valid;
output 	src_payload;
output 	src_payload1;
output 	src_payload2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \saved_grant[1]~0_combout ;


dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\saved_grant[1]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cyclonev_lcell_comb \src_valid~0 (
	.dataa(!h2f_ARVALID_0),
	.datab(!has_pending_responses),
	.datac(!saved_grant_1),
	.datad(!Equal7),
	.datae(!last_channel_7),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~0 .extended_lut = "off";
defparam \src_valid~0 .lut_mask = 64'h0004000500040005;
defparam \src_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!h2f_ARSIZE_0),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h1111111111111111;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!h2f_ARSIZE_1),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h1111111111111111;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!h2f_ARSIZE_2),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h1111111111111111;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!nxt_in_ready),
	.datab(!\packet_in_progress~q ),
	.datac(!src_valid),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'h3535353535353535;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \saved_grant[1]~0 (
	.dataa(!h2f_ARVALID_0),
	.datab(!has_pending_responses),
	.datac(!saved_grant_1),
	.datad(!Equal7),
	.datae(!last_channel_7),
	.dataf(!\packet_in_progress~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\saved_grant[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \saved_grant[1]~0 .extended_lut = "off";
defparam \saved_grant[1]~0 .lut_mask = 64'h004400550F0F0F0F;
defparam \saved_grant[1]~0 .shared_arith = "off";

endmodule

module spw_babasu_spw_babasu_mm_interconnect_0_cmd_mux_8 (
	h2f_ARVALID_0,
	h2f_ARSIZE_0,
	h2f_ARSIZE_1,
	h2f_ARSIZE_2,
	has_pending_responses,
	saved_grant_1,
	src_channel,
	altera_reset_synchronizer_int_chain_out,
	nxt_in_ready,
	last_channel_8,
	src_valid,
	src_payload,
	src_payload1,
	src_payload2,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARVALID_0;
input 	h2f_ARSIZE_0;
input 	h2f_ARSIZE_1;
input 	h2f_ARSIZE_2;
input 	has_pending_responses;
output 	saved_grant_1;
input 	src_channel;
input 	altera_reset_synchronizer_int_chain_out;
input 	nxt_in_ready;
input 	last_channel_8;
output 	src_valid;
output 	src_payload;
output 	src_payload1;
output 	src_payload2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \saved_grant[1]~0_combout ;
wire \saved_grant[1]~1_combout ;


dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\saved_grant[1]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cyclonev_lcell_comb \src_valid~0 (
	.dataa(!saved_grant_1),
	.datab(!src_channel),
	.datac(!\saved_grant[1]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~0 .extended_lut = "off";
defparam \src_valid~0 .lut_mask = 64'h0101010101010101;
defparam \src_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!h2f_ARSIZE_0),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h1111111111111111;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!h2f_ARSIZE_2),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h1111111111111111;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!h2f_ARSIZE_1),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h1111111111111111;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!nxt_in_ready),
	.datab(!\packet_in_progress~q ),
	.datac(!src_valid),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'h3535353535353535;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \saved_grant[1]~0 (
	.dataa(!h2f_ARVALID_0),
	.datab(!has_pending_responses),
	.datac(!last_channel_8),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\saved_grant[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \saved_grant[1]~0 .extended_lut = "off";
defparam \saved_grant[1]~0 .lut_mask = 64'h4545454545454545;
defparam \saved_grant[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \saved_grant[1]~1 (
	.dataa(!saved_grant_1),
	.datab(!src_channel),
	.datac(gnd),
	.datad(!\packet_in_progress~q ),
	.datae(!\saved_grant[1]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\saved_grant[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \saved_grant[1]~1 .extended_lut = "off";
defparam \saved_grant[1]~1 .lut_mask = 64'h0055335500553355;
defparam \saved_grant[1]~1 .shared_arith = "off";

endmodule

module spw_babasu_spw_babasu_mm_interconnect_0_cmd_mux_9 (
	h2f_WLAST_0,
	h2f_ARID_0,
	h2f_ARID_1,
	h2f_ARID_2,
	h2f_ARID_3,
	h2f_ARID_4,
	h2f_ARID_5,
	h2f_ARID_6,
	h2f_ARID_7,
	h2f_ARID_8,
	h2f_ARID_9,
	h2f_ARID_10,
	h2f_ARID_11,
	h2f_ARSIZE_0,
	h2f_ARSIZE_1,
	h2f_ARSIZE_2,
	h2f_AWID_0,
	h2f_AWID_1,
	h2f_AWID_2,
	h2f_AWID_3,
	h2f_AWID_4,
	h2f_AWID_5,
	h2f_AWID_6,
	h2f_AWID_7,
	h2f_AWID_8,
	h2f_AWID_9,
	h2f_AWID_10,
	h2f_AWID_11,
	h2f_AWSIZE_0,
	h2f_AWSIZE_1,
	h2f_AWSIZE_2,
	h2f_WDATA_0,
	h2f_WSTRB_0,
	h2f_WSTRB_1,
	h2f_WSTRB_2,
	h2f_WSTRB_3,
	nxt_in_ready,
	nxt_in_ready1,
	saved_grant_1,
	write_addr_data_both_valid,
	out_data_5,
	Equal15,
	Equal9,
	saved_grant_0,
	altera_reset_synchronizer_int_chain_out,
	Equal5,
	src9_valid,
	src9_valid1,
	Equal91,
	src9_valid2,
	src_valid,
	src_data_87,
	src_data_88,
	src_valid1,
	src_data_35,
	src_data_34,
	src_data_33,
	src_data_32,
	src_payload_0,
	src9_valid3,
	src9_valid4,
	Selector3,
	Selector10,
	Selector4,
	Selector11,
	src_payload,
	src_data_82,
	src_data_81,
	src_data_105,
	src_data_106,
	src_data_107,
	src_data_108,
	src_data_109,
	src_data_110,
	src_data_111,
	src_data_112,
	src_data_113,
	src_data_114,
	src_data_115,
	src_data_116,
	src_data_86,
	Selector5,
	Selector12,
	src_data_80,
	Selector6,
	Selector13,
	src_data_79,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_WLAST_0;
input 	h2f_ARID_0;
input 	h2f_ARID_1;
input 	h2f_ARID_2;
input 	h2f_ARID_3;
input 	h2f_ARID_4;
input 	h2f_ARID_5;
input 	h2f_ARID_6;
input 	h2f_ARID_7;
input 	h2f_ARID_8;
input 	h2f_ARID_9;
input 	h2f_ARID_10;
input 	h2f_ARID_11;
input 	h2f_ARSIZE_0;
input 	h2f_ARSIZE_1;
input 	h2f_ARSIZE_2;
input 	h2f_AWID_0;
input 	h2f_AWID_1;
input 	h2f_AWID_2;
input 	h2f_AWID_3;
input 	h2f_AWID_4;
input 	h2f_AWID_5;
input 	h2f_AWID_6;
input 	h2f_AWID_7;
input 	h2f_AWID_8;
input 	h2f_AWID_9;
input 	h2f_AWID_10;
input 	h2f_AWID_11;
input 	h2f_AWSIZE_0;
input 	h2f_AWSIZE_1;
input 	h2f_AWSIZE_2;
input 	h2f_WDATA_0;
input 	h2f_WSTRB_0;
input 	h2f_WSTRB_1;
input 	h2f_WSTRB_2;
input 	h2f_WSTRB_3;
input 	nxt_in_ready;
input 	nxt_in_ready1;
output 	saved_grant_1;
input 	write_addr_data_both_valid;
input 	out_data_5;
input 	Equal15;
input 	Equal9;
output 	saved_grant_0;
input 	altera_reset_synchronizer_int_chain_out;
input 	Equal5;
input 	src9_valid;
input 	src9_valid1;
input 	Equal91;
input 	src9_valid2;
output 	src_valid;
output 	src_data_87;
output 	src_data_88;
output 	src_valid1;
output 	src_data_35;
output 	src_data_34;
output 	src_data_33;
output 	src_data_32;
output 	src_payload_0;
input 	src9_valid3;
input 	src9_valid4;
input 	Selector3;
input 	Selector10;
input 	Selector4;
input 	Selector11;
output 	src_payload;
output 	src_data_82;
output 	src_data_81;
output 	src_data_105;
output 	src_data_106;
output 	src_data_107;
output 	src_data_108;
output 	src_data_109;
output 	src_data_110;
output 	src_data_111;
output 	src_data_112;
output 	src_data_113;
output 	src_data_114;
output 	src_data_115;
output 	src_data_116;
output 	src_data_86;
input 	Selector5;
input 	Selector12;
output 	src_data_80;
input 	Selector6;
input 	Selector13;
output 	src_data_79;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[1]~0_combout ;
wire \arb|grant[0]~1_combout ;
wire \WideOr1~combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~0_combout ;


spw_babasu_altera_merlin_arbitrator_8 arb(
	.nxt_in_ready(nxt_in_ready),
	.nxt_in_ready1(nxt_in_ready1),
	.Equal9(Equal9),
	.reset(altera_reset_synchronizer_int_chain_out),
	.Equal5(Equal5),
	.src9_valid(src9_valid1),
	.src_payload_0(src_payload_0),
	.src9_valid1(src9_valid3),
	.src9_valid2(src9_valid4),
	.grant_1(\arb|grant[1]~0_combout ),
	.packet_in_progress(\packet_in_progress~q ),
	.grant_0(\arb|grant[0]~1_combout ),
	.WideOr1(\WideOr1~combout ),
	.clk(clk_clk));

cyclonev_lcell_comb WideOr1(
	.dataa(!Equal5),
	.datab(!Equal9),
	.datac(!saved_grant_0),
	.datad(!src9_valid1),
	.datae(!src_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr1.extended_lut = "off";
defparam WideOr1.lut_mask = 64'hFFFE0000FFFE0000;
defparam WideOr1.shared_arith = "off";

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

cyclonev_lcell_comb \src_valid~0 (
	.dataa(!saved_grant_1),
	.datab(!Equal91),
	.datac(!src9_valid2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~0 .extended_lut = "off";
defparam \src_valid~0 .lut_mask = 64'h0101010101010101;
defparam \src_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[87] (
	.dataa(!h2f_ARSIZE_1),
	.datab(!h2f_AWSIZE_1),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_87),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[87] .extended_lut = "off";
defparam \src_data[87] .lut_mask = 64'h0537053705370537;
defparam \src_data[87] .shared_arith = "off";

cyclonev_lcell_comb \src_data[88] (
	.dataa(!h2f_ARSIZE_2),
	.datab(!h2f_AWSIZE_2),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_88),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[88] .extended_lut = "off";
defparam \src_data[88] .lut_mask = 64'h0537053705370537;
defparam \src_data[88] .shared_arith = "off";

cyclonev_lcell_comb \src_valid~1 (
	.dataa(!out_data_5),
	.datab(!Equal15),
	.datac(!Equal9),
	.datad(!saved_grant_0),
	.datae(!write_addr_data_both_valid),
	.dataf(!src9_valid),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~1 .extended_lut = "off";
defparam \src_valid~1 .lut_mask = 64'h0000000200000000;
defparam \src_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \src_data[35] (
	.dataa(!h2f_WSTRB_3),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_35),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[35] .extended_lut = "off";
defparam \src_data[35] .lut_mask = 64'h3737373737373737;
defparam \src_data[35] .shared_arith = "off";

cyclonev_lcell_comb \src_data[34] (
	.dataa(!h2f_WSTRB_2),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_34),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[34] .extended_lut = "off";
defparam \src_data[34] .lut_mask = 64'h3737373737373737;
defparam \src_data[34] .shared_arith = "off";

cyclonev_lcell_comb \src_data[33] (
	.dataa(!h2f_WSTRB_1),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_33),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[33] .extended_lut = "off";
defparam \src_data[33] .lut_mask = 64'h3737373737373737;
defparam \src_data[33] .shared_arith = "off";

cyclonev_lcell_comb \src_data[32] (
	.dataa(!h2f_WSTRB_0),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_32),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[32] .extended_lut = "off";
defparam \src_data[32] .lut_mask = 64'h3737373737373737;
defparam \src_data[32] .shared_arith = "off";

cyclonev_lcell_comb \src_payload[0] (
	.dataa(!h2f_WLAST_0),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload[0] .extended_lut = "off";
defparam \src_payload[0] .lut_mask = 64'h3737373737373737;
defparam \src_payload[0] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!h2f_WDATA_0),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h1111111111111111;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[82] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector3),
	.datad(!Selector10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_82),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[82] .extended_lut = "off";
defparam \src_data[82] .lut_mask = 64'h0357035703570357;
defparam \src_data[82] .shared_arith = "off";

cyclonev_lcell_comb \src_data[81] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector4),
	.datad(!Selector11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_81),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[81] .extended_lut = "off";
defparam \src_data[81] .lut_mask = 64'h0357035703570357;
defparam \src_data[81] .shared_arith = "off";

cyclonev_lcell_comb \src_data[105] (
	.dataa(!h2f_ARID_0),
	.datab(!h2f_AWID_0),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_105),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[105] .extended_lut = "off";
defparam \src_data[105] .lut_mask = 64'h0537053705370537;
defparam \src_data[105] .shared_arith = "off";

cyclonev_lcell_comb \src_data[106] (
	.dataa(!h2f_ARID_1),
	.datab(!h2f_AWID_1),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_106),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[106] .extended_lut = "off";
defparam \src_data[106] .lut_mask = 64'h0537053705370537;
defparam \src_data[106] .shared_arith = "off";

cyclonev_lcell_comb \src_data[107] (
	.dataa(!h2f_ARID_2),
	.datab(!h2f_AWID_2),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_107),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[107] .extended_lut = "off";
defparam \src_data[107] .lut_mask = 64'h0537053705370537;
defparam \src_data[107] .shared_arith = "off";

cyclonev_lcell_comb \src_data[108] (
	.dataa(!h2f_ARID_3),
	.datab(!h2f_AWID_3),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_108),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[108] .extended_lut = "off";
defparam \src_data[108] .lut_mask = 64'h0537053705370537;
defparam \src_data[108] .shared_arith = "off";

cyclonev_lcell_comb \src_data[109] (
	.dataa(!h2f_ARID_4),
	.datab(!h2f_AWID_4),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_109),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[109] .extended_lut = "off";
defparam \src_data[109] .lut_mask = 64'h0537053705370537;
defparam \src_data[109] .shared_arith = "off";

cyclonev_lcell_comb \src_data[110] (
	.dataa(!h2f_ARID_5),
	.datab(!h2f_AWID_5),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_110),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[110] .extended_lut = "off";
defparam \src_data[110] .lut_mask = 64'h0537053705370537;
defparam \src_data[110] .shared_arith = "off";

cyclonev_lcell_comb \src_data[111] (
	.dataa(!h2f_ARID_6),
	.datab(!h2f_AWID_6),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_111),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[111] .extended_lut = "off";
defparam \src_data[111] .lut_mask = 64'h0537053705370537;
defparam \src_data[111] .shared_arith = "off";

cyclonev_lcell_comb \src_data[112] (
	.dataa(!h2f_ARID_7),
	.datab(!h2f_AWID_7),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_112),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[112] .extended_lut = "off";
defparam \src_data[112] .lut_mask = 64'h0537053705370537;
defparam \src_data[112] .shared_arith = "off";

cyclonev_lcell_comb \src_data[113] (
	.dataa(!h2f_ARID_8),
	.datab(!h2f_AWID_8),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_113),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[113] .extended_lut = "off";
defparam \src_data[113] .lut_mask = 64'h0537053705370537;
defparam \src_data[113] .shared_arith = "off";

cyclonev_lcell_comb \src_data[114] (
	.dataa(!h2f_ARID_9),
	.datab(!h2f_AWID_9),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_114),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[114] .extended_lut = "off";
defparam \src_data[114] .lut_mask = 64'h0537053705370537;
defparam \src_data[114] .shared_arith = "off";

cyclonev_lcell_comb \src_data[115] (
	.dataa(!h2f_ARID_10),
	.datab(!h2f_AWID_10),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_115),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[115] .extended_lut = "off";
defparam \src_data[115] .lut_mask = 64'h0537053705370537;
defparam \src_data[115] .shared_arith = "off";

cyclonev_lcell_comb \src_data[116] (
	.dataa(!h2f_ARID_11),
	.datab(!h2f_AWID_11),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_116),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[116] .extended_lut = "off";
defparam \src_data[116] .lut_mask = 64'h0537053705370537;
defparam \src_data[116] .shared_arith = "off";

cyclonev_lcell_comb \src_data[86] (
	.dataa(!h2f_ARSIZE_0),
	.datab(!h2f_AWSIZE_0),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_86),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[86] .extended_lut = "off";
defparam \src_data[86] .lut_mask = 64'h0537053705370537;
defparam \src_data[86] .shared_arith = "off";

cyclonev_lcell_comb \src_data[80] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector5),
	.datad(!Selector12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_80),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[80] .extended_lut = "off";
defparam \src_data[80] .lut_mask = 64'h0357035703570357;
defparam \src_data[80] .shared_arith = "off";

cyclonev_lcell_comb \src_data[79] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector6),
	.datad(!Selector13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_79),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[79] .extended_lut = "off";
defparam \src_data[79] .lut_mask = 64'h0357035703570357;
defparam \src_data[79] .shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!\update_grant~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \update_grant~0 (
	.dataa(!nxt_in_ready1),
	.datab(!nxt_in_ready),
	.datac(!src_valid),
	.datad(!src_valid1),
	.datae(!src_payload_0),
	.dataf(!\packet_in_progress~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\update_grant~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \update_grant~0 .extended_lut = "off";
defparam \update_grant~0 .lut_mask = 64'hF000F77700000777;
defparam \update_grant~0 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_arbitrator_8 (
	nxt_in_ready,
	nxt_in_ready1,
	Equal9,
	reset,
	Equal5,
	src9_valid,
	src_payload_0,
	src9_valid1,
	src9_valid2,
	grant_1,
	packet_in_progress,
	grant_0,
	WideOr1,
	clk)/* synthesis synthesis_greybox=0 */;
input 	nxt_in_ready;
input 	nxt_in_ready1;
input 	Equal9;
input 	reset;
input 	Equal5;
input 	src9_valid;
input 	src_payload_0;
input 	src9_valid1;
input 	src9_valid2;
output 	grant_1;
input 	packet_in_progress;
output 	grant_0;
input 	WideOr1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg[0]~2_combout ;
wire \top_priority_reg[0]~q ;


cyclonev_lcell_comb \grant[1]~0 (
	.dataa(!\top_priority_reg[1]~q ),
	.datab(!\top_priority_reg[0]~q ),
	.datac(!src9_valid1),
	.datad(!src9_valid2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[1]~0 .extended_lut = "off";
defparam \grant[1]~0 .lut_mask = 64'h00D500D500D500D5;
defparam \grant[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \grant[0]~1 (
	.dataa(!\top_priority_reg[1]~q ),
	.datab(!\top_priority_reg[0]~q ),
	.datac(!src9_valid1),
	.datad(!src9_valid2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[0]~1 .extended_lut = "off";
defparam \grant[0]~1 .lut_mask = 64'h0D0C0D0C0D0C0D0C;
defparam \grant[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~0 (
	.dataa(!Equal5),
	.datab(!Equal9),
	.datac(!src9_valid),
	.datad(!src9_valid2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~0 .extended_lut = "off";
defparam \top_priority_reg[0]~0 .lut_mask = 64'hFE00FE00FE00FE00;
defparam \top_priority_reg[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~1 (
	.dataa(!nxt_in_ready1),
	.datab(!nxt_in_ready),
	.datac(!WideOr1),
	.datad(!src_payload_0),
	.datae(!packet_in_progress),
	.dataf(!\top_priority_reg[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~1 .extended_lut = "off";
defparam \top_priority_reg[0]~1 .lut_mask = 64'h0F7F007000000000;
defparam \top_priority_reg[0]~1 .shared_arith = "off";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~1_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

cyclonev_lcell_comb \top_priority_reg[0]~2 (
	.dataa(!grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~2 .extended_lut = "off";
defparam \top_priority_reg[0]~2 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \top_priority_reg[0]~2 .shared_arith = "off";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~1_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

endmodule

module spw_babasu_spw_babasu_mm_interconnect_0_cmd_mux_10 (
	h2f_ARVALID_0,
	h2f_ARSIZE_0,
	h2f_ARSIZE_1,
	h2f_ARSIZE_2,
	has_pending_responses,
	saved_grant_1,
	Equal10,
	altera_reset_synchronizer_int_chain_out,
	last_channel_10,
	src_valid,
	nxt_in_ready,
	src_payload,
	src_payload1,
	src_payload2,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARVALID_0;
input 	h2f_ARSIZE_0;
input 	h2f_ARSIZE_1;
input 	h2f_ARSIZE_2;
input 	has_pending_responses;
output 	saved_grant_1;
input 	Equal10;
input 	altera_reset_synchronizer_int_chain_out;
input 	last_channel_10;
output 	src_valid;
input 	nxt_in_ready;
output 	src_payload;
output 	src_payload1;
output 	src_payload2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \saved_grant[1]~0_combout ;


dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\saved_grant[1]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cyclonev_lcell_comb \src_valid~0 (
	.dataa(!h2f_ARVALID_0),
	.datab(!has_pending_responses),
	.datac(!saved_grant_1),
	.datad(!Equal10),
	.datae(!last_channel_10),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~0 .extended_lut = "off";
defparam \src_valid~0 .lut_mask = 64'h0004000500040005;
defparam \src_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!h2f_ARSIZE_0),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h1111111111111111;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!h2f_ARSIZE_1),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h1111111111111111;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!h2f_ARSIZE_2),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h1111111111111111;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!nxt_in_ready),
	.datab(!\packet_in_progress~q ),
	.datac(!src_valid),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'h3535353535353535;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \saved_grant[1]~0 (
	.dataa(!h2f_ARVALID_0),
	.datab(!has_pending_responses),
	.datac(!saved_grant_1),
	.datad(!Equal10),
	.datae(!last_channel_10),
	.dataf(!\packet_in_progress~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\saved_grant[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \saved_grant[1]~0 .extended_lut = "off";
defparam \saved_grant[1]~0 .lut_mask = 64'h004400550F0F0F0F;
defparam \saved_grant[1]~0 .shared_arith = "off";

endmodule

module spw_babasu_spw_babasu_mm_interconnect_0_cmd_mux_11 (
	h2f_ARVALID_0,
	h2f_ARADDR_4,
	h2f_ARADDR_5,
	h2f_ARADDR_6,
	h2f_ARADDR_7,
	h2f_ARADDR_8,
	h2f_ARSIZE_0,
	h2f_ARSIZE_1,
	h2f_ARSIZE_2,
	has_pending_responses,
	saved_grant_1,
	last_cycle,
	altera_reset_synchronizer_int_chain_out,
	nxt_in_ready,
	last_channel_11,
	src_valid,
	src_payload,
	src_payload1,
	src_payload2,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARVALID_0;
input 	h2f_ARADDR_4;
input 	h2f_ARADDR_5;
input 	h2f_ARADDR_6;
input 	h2f_ARADDR_7;
input 	h2f_ARADDR_8;
input 	h2f_ARSIZE_0;
input 	h2f_ARSIZE_1;
input 	h2f_ARSIZE_2;
input 	has_pending_responses;
output 	saved_grant_1;
output 	last_cycle;
input 	altera_reset_synchronizer_int_chain_out;
input 	nxt_in_ready;
input 	last_channel_11;
output 	src_valid;
output 	src_payload;
output 	src_payload1;
output 	src_payload2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \saved_grant[1]~0_combout ;
wire \saved_grant[1]~1_combout ;


dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\saved_grant[1]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cyclonev_lcell_comb \last_cycle~0 (
	.dataa(!h2f_ARADDR_4),
	.datab(!h2f_ARADDR_5),
	.datac(!h2f_ARADDR_6),
	.datad(!h2f_ARADDR_7),
	.datae(!h2f_ARADDR_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_cycle),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_cycle~0 .extended_lut = "off";
defparam \last_cycle~0 .lut_mask = 64'h0010000000100000;
defparam \last_cycle~0 .shared_arith = "off";

cyclonev_lcell_comb \src_valid~0 (
	.dataa(!saved_grant_1),
	.datab(!last_cycle),
	.datac(!\saved_grant[1]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~0 .extended_lut = "off";
defparam \src_valid~0 .lut_mask = 64'h0101010101010101;
defparam \src_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!h2f_ARSIZE_0),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h1111111111111111;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!h2f_ARSIZE_2),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h1111111111111111;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!h2f_ARSIZE_1),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h1111111111111111;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!nxt_in_ready),
	.datab(!\packet_in_progress~q ),
	.datac(!src_valid),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'h3535353535353535;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \saved_grant[1]~0 (
	.dataa(!h2f_ARVALID_0),
	.datab(!has_pending_responses),
	.datac(!last_channel_11),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\saved_grant[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \saved_grant[1]~0 .extended_lut = "off";
defparam \saved_grant[1]~0 .lut_mask = 64'h4545454545454545;
defparam \saved_grant[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \saved_grant[1]~1 (
	.dataa(!saved_grant_1),
	.datab(!last_cycle),
	.datac(gnd),
	.datad(!\packet_in_progress~q ),
	.datae(!\saved_grant[1]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\saved_grant[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \saved_grant[1]~1 .extended_lut = "off";
defparam \saved_grant[1]~1 .lut_mask = 64'h0055335500553355;
defparam \saved_grant[1]~1 .shared_arith = "off";

endmodule

module spw_babasu_spw_babasu_mm_interconnect_0_cmd_mux_12 (
	h2f_ARVALID_0,
	h2f_ARADDR_4,
	h2f_ARADDR_5,
	h2f_ARADDR_6,
	h2f_ARADDR_7,
	h2f_ARADDR_8,
	h2f_ARSIZE_0,
	h2f_ARSIZE_1,
	h2f_ARSIZE_2,
	has_pending_responses,
	saved_grant_1,
	last_cycle,
	altera_reset_synchronizer_int_chain_out,
	nxt_in_ready,
	last_channel_12,
	src_valid,
	src_payload,
	src_payload1,
	src_payload2,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARVALID_0;
input 	h2f_ARADDR_4;
input 	h2f_ARADDR_5;
input 	h2f_ARADDR_6;
input 	h2f_ARADDR_7;
input 	h2f_ARADDR_8;
input 	h2f_ARSIZE_0;
input 	h2f_ARSIZE_1;
input 	h2f_ARSIZE_2;
input 	has_pending_responses;
output 	saved_grant_1;
output 	last_cycle;
input 	altera_reset_synchronizer_int_chain_out;
input 	nxt_in_ready;
input 	last_channel_12;
output 	src_valid;
output 	src_payload;
output 	src_payload1;
output 	src_payload2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \saved_grant[1]~0_combout ;
wire \saved_grant[1]~1_combout ;


dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\saved_grant[1]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cyclonev_lcell_comb \last_cycle~0 (
	.dataa(!h2f_ARADDR_4),
	.datab(!h2f_ARADDR_5),
	.datac(!h2f_ARADDR_6),
	.datad(!h2f_ARADDR_7),
	.datae(!h2f_ARADDR_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_cycle),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_cycle~0 .extended_lut = "off";
defparam \last_cycle~0 .lut_mask = 64'h0008000000080000;
defparam \last_cycle~0 .shared_arith = "off";

cyclonev_lcell_comb \src_valid~0 (
	.dataa(!saved_grant_1),
	.datab(!last_cycle),
	.datac(!\saved_grant[1]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~0 .extended_lut = "off";
defparam \src_valid~0 .lut_mask = 64'h0101010101010101;
defparam \src_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!h2f_ARSIZE_0),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h1111111111111111;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!h2f_ARSIZE_1),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h1111111111111111;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!h2f_ARSIZE_2),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h1111111111111111;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!nxt_in_ready),
	.datab(!\packet_in_progress~q ),
	.datac(!src_valid),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'h3535353535353535;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \saved_grant[1]~0 (
	.dataa(!h2f_ARVALID_0),
	.datab(!has_pending_responses),
	.datac(!last_channel_12),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\saved_grant[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \saved_grant[1]~0 .extended_lut = "off";
defparam \saved_grant[1]~0 .lut_mask = 64'h4545454545454545;
defparam \saved_grant[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \saved_grant[1]~1 (
	.dataa(!saved_grant_1),
	.datab(!last_cycle),
	.datac(gnd),
	.datad(!\packet_in_progress~q ),
	.datae(!\saved_grant[1]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\saved_grant[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \saved_grant[1]~1 .extended_lut = "off";
defparam \saved_grant[1]~1 .lut_mask = 64'h0055335500553355;
defparam \saved_grant[1]~1 .shared_arith = "off";

endmodule

module spw_babasu_spw_babasu_mm_interconnect_0_cmd_mux_13 (
	h2f_ARVALID_0,
	h2f_WLAST_0,
	h2f_ARADDR_4,
	h2f_ARADDR_5,
	h2f_ARADDR_6,
	h2f_ARADDR_7,
	h2f_ARADDR_8,
	h2f_ARID_0,
	h2f_ARID_1,
	h2f_ARID_2,
	h2f_ARID_3,
	h2f_ARID_4,
	h2f_ARID_5,
	h2f_ARID_6,
	h2f_ARID_7,
	h2f_ARID_8,
	h2f_ARID_9,
	h2f_ARID_10,
	h2f_ARID_11,
	h2f_ARSIZE_0,
	h2f_ARSIZE_1,
	h2f_ARSIZE_2,
	h2f_AWID_0,
	h2f_AWID_1,
	h2f_AWID_2,
	h2f_AWID_3,
	h2f_AWID_4,
	h2f_AWID_5,
	h2f_AWID_6,
	h2f_AWID_7,
	h2f_AWID_8,
	h2f_AWID_9,
	h2f_AWID_10,
	h2f_AWID_11,
	h2f_AWSIZE_0,
	h2f_AWSIZE_1,
	h2f_AWSIZE_2,
	h2f_WDATA_0,
	h2f_WSTRB_0,
	h2f_WSTRB_1,
	h2f_WSTRB_2,
	h2f_WSTRB_3,
	nxt_in_ready,
	has_pending_responses,
	nxt_in_ready1,
	saved_grant_1,
	write_addr_data_both_valid,
	out_data_5,
	Equal13,
	Equal15,
	saved_grant_0,
	altera_reset_synchronizer_int_chain_out,
	Equal5,
	src13_valid,
	src13_valid1,
	last_channel_13,
	src_valid,
	src_data_87,
	src_data_88,
	src_valid1,
	src_data_35,
	src_data_34,
	src_data_33,
	src_data_32,
	src_payload_0,
	src13_valid2,
	Selector3,
	Selector10,
	Selector4,
	Selector11,
	src_payload,
	src_data_82,
	src_data_81,
	src_data_105,
	src_data_106,
	src_data_107,
	src_data_108,
	src_data_109,
	src_data_110,
	src_data_111,
	src_data_112,
	src_data_113,
	src_data_114,
	src_data_115,
	src_data_116,
	src_data_86,
	Selector5,
	Selector12,
	src_data_80,
	Selector6,
	Selector13,
	src_data_79,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARVALID_0;
input 	h2f_WLAST_0;
input 	h2f_ARADDR_4;
input 	h2f_ARADDR_5;
input 	h2f_ARADDR_6;
input 	h2f_ARADDR_7;
input 	h2f_ARADDR_8;
input 	h2f_ARID_0;
input 	h2f_ARID_1;
input 	h2f_ARID_2;
input 	h2f_ARID_3;
input 	h2f_ARID_4;
input 	h2f_ARID_5;
input 	h2f_ARID_6;
input 	h2f_ARID_7;
input 	h2f_ARID_8;
input 	h2f_ARID_9;
input 	h2f_ARID_10;
input 	h2f_ARID_11;
input 	h2f_ARSIZE_0;
input 	h2f_ARSIZE_1;
input 	h2f_ARSIZE_2;
input 	h2f_AWID_0;
input 	h2f_AWID_1;
input 	h2f_AWID_2;
input 	h2f_AWID_3;
input 	h2f_AWID_4;
input 	h2f_AWID_5;
input 	h2f_AWID_6;
input 	h2f_AWID_7;
input 	h2f_AWID_8;
input 	h2f_AWID_9;
input 	h2f_AWID_10;
input 	h2f_AWID_11;
input 	h2f_AWSIZE_0;
input 	h2f_AWSIZE_1;
input 	h2f_AWSIZE_2;
input 	h2f_WDATA_0;
input 	h2f_WSTRB_0;
input 	h2f_WSTRB_1;
input 	h2f_WSTRB_2;
input 	h2f_WSTRB_3;
input 	nxt_in_ready;
input 	has_pending_responses;
input 	nxt_in_ready1;
output 	saved_grant_1;
input 	write_addr_data_both_valid;
input 	out_data_5;
input 	Equal13;
input 	Equal15;
output 	saved_grant_0;
input 	altera_reset_synchronizer_int_chain_out;
input 	Equal5;
input 	src13_valid;
input 	src13_valid1;
input 	last_channel_13;
output 	src_valid;
output 	src_data_87;
output 	src_data_88;
output 	src_valid1;
output 	src_data_35;
output 	src_data_34;
output 	src_data_33;
output 	src_data_32;
output 	src_payload_0;
input 	src13_valid2;
input 	Selector3;
input 	Selector10;
input 	Selector4;
input 	Selector11;
output 	src_payload;
output 	src_data_82;
output 	src_data_81;
output 	src_data_105;
output 	src_data_106;
output 	src_data_107;
output 	src_data_108;
output 	src_data_109;
output 	src_data_110;
output 	src_data_111;
output 	src_data_112;
output 	src_data_113;
output 	src_data_114;
output 	src_data_115;
output 	src_data_116;
output 	src_data_86;
input 	Selector5;
input 	Selector12;
output 	src_data_80;
input 	Selector6;
input 	Selector13;
output 	src_data_79;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \src_valid~4_combout ;
wire \arb|grant[1]~0_combout ;
wire \arb|grant[0]~1_combout ;
wire \WideOr1~combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~0_combout ;
wire \src_valid~0_combout ;
wire \src_valid~1_combout ;


spw_babasu_altera_merlin_arbitrator_12 arb(
	.nxt_in_ready(nxt_in_ready),
	.nxt_in_ready1(nxt_in_ready1),
	.Equal13(Equal13),
	.reset(altera_reset_synchronizer_int_chain_out),
	.Equal5(Equal5),
	.src13_valid(src13_valid1),
	.src_payload_0(src_payload_0),
	.src13_valid1(src13_valid2),
	.src_valid(\src_valid~4_combout ),
	.grant_1(\arb|grant[1]~0_combout ),
	.packet_in_progress(\packet_in_progress~q ),
	.grant_0(\arb|grant[0]~1_combout ),
	.WideOr1(\WideOr1~combout ),
	.clk(clk_clk));

cyclonev_lcell_comb \src_valid~4 (
	.dataa(!\src_valid~0_combout ),
	.datab(!\src_valid~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_valid~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~4 .extended_lut = "off";
defparam \src_valid~4 .lut_mask = 64'h1111111111111111;
defparam \src_valid~4 .shared_arith = "off";

cyclonev_lcell_comb WideOr1(
	.dataa(!Equal5),
	.datab(!Equal13),
	.datac(!saved_grant_0),
	.datad(!src13_valid1),
	.datae(!src_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr1.extended_lut = "off";
defparam WideOr1.lut_mask = 64'hFFFE0000FFFE0000;
defparam WideOr1.shared_arith = "off";

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

cyclonev_lcell_comb \src_valid~2 (
	.dataa(!saved_grant_1),
	.datab(!\src_valid~0_combout ),
	.datac(!\src_valid~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~2 .extended_lut = "off";
defparam \src_valid~2 .lut_mask = 64'h0101010101010101;
defparam \src_valid~2 .shared_arith = "off";

cyclonev_lcell_comb \src_data[87] (
	.dataa(!h2f_ARSIZE_1),
	.datab(!h2f_AWSIZE_1),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_87),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[87] .extended_lut = "off";
defparam \src_data[87] .lut_mask = 64'h0537053705370537;
defparam \src_data[87] .shared_arith = "off";

cyclonev_lcell_comb \src_data[88] (
	.dataa(!h2f_ARSIZE_2),
	.datab(!h2f_AWSIZE_2),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_88),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[88] .extended_lut = "off";
defparam \src_data[88] .lut_mask = 64'h0537053705370537;
defparam \src_data[88] .shared_arith = "off";

cyclonev_lcell_comb \src_valid~3 (
	.dataa(!out_data_5),
	.datab(!Equal15),
	.datac(!Equal13),
	.datad(!saved_grant_0),
	.datae(!write_addr_data_both_valid),
	.dataf(!src13_valid),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~3 .extended_lut = "off";
defparam \src_valid~3 .lut_mask = 64'h0000000200000000;
defparam \src_valid~3 .shared_arith = "off";

cyclonev_lcell_comb \src_data[35] (
	.dataa(!h2f_WSTRB_3),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_35),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[35] .extended_lut = "off";
defparam \src_data[35] .lut_mask = 64'h3737373737373737;
defparam \src_data[35] .shared_arith = "off";

cyclonev_lcell_comb \src_data[34] (
	.dataa(!h2f_WSTRB_2),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_34),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[34] .extended_lut = "off";
defparam \src_data[34] .lut_mask = 64'h3737373737373737;
defparam \src_data[34] .shared_arith = "off";

cyclonev_lcell_comb \src_data[33] (
	.dataa(!h2f_WSTRB_1),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_33),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[33] .extended_lut = "off";
defparam \src_data[33] .lut_mask = 64'h3737373737373737;
defparam \src_data[33] .shared_arith = "off";

cyclonev_lcell_comb \src_data[32] (
	.dataa(!h2f_WSTRB_0),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_32),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[32] .extended_lut = "off";
defparam \src_data[32] .lut_mask = 64'h3737373737373737;
defparam \src_data[32] .shared_arith = "off";

cyclonev_lcell_comb \src_payload[0] (
	.dataa(!h2f_WLAST_0),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload[0] .extended_lut = "off";
defparam \src_payload[0] .lut_mask = 64'h3737373737373737;
defparam \src_payload[0] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!h2f_WDATA_0),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h1111111111111111;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[82] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector3),
	.datad(!Selector10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_82),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[82] .extended_lut = "off";
defparam \src_data[82] .lut_mask = 64'h0357035703570357;
defparam \src_data[82] .shared_arith = "off";

cyclonev_lcell_comb \src_data[81] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector4),
	.datad(!Selector11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_81),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[81] .extended_lut = "off";
defparam \src_data[81] .lut_mask = 64'h0357035703570357;
defparam \src_data[81] .shared_arith = "off";

cyclonev_lcell_comb \src_data[105] (
	.dataa(!h2f_ARID_0),
	.datab(!h2f_AWID_0),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_105),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[105] .extended_lut = "off";
defparam \src_data[105] .lut_mask = 64'h0537053705370537;
defparam \src_data[105] .shared_arith = "off";

cyclonev_lcell_comb \src_data[106] (
	.dataa(!h2f_ARID_1),
	.datab(!h2f_AWID_1),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_106),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[106] .extended_lut = "off";
defparam \src_data[106] .lut_mask = 64'h0537053705370537;
defparam \src_data[106] .shared_arith = "off";

cyclonev_lcell_comb \src_data[107] (
	.dataa(!h2f_ARID_2),
	.datab(!h2f_AWID_2),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_107),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[107] .extended_lut = "off";
defparam \src_data[107] .lut_mask = 64'h0537053705370537;
defparam \src_data[107] .shared_arith = "off";

cyclonev_lcell_comb \src_data[108] (
	.dataa(!h2f_ARID_3),
	.datab(!h2f_AWID_3),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_108),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[108] .extended_lut = "off";
defparam \src_data[108] .lut_mask = 64'h0537053705370537;
defparam \src_data[108] .shared_arith = "off";

cyclonev_lcell_comb \src_data[109] (
	.dataa(!h2f_ARID_4),
	.datab(!h2f_AWID_4),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_109),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[109] .extended_lut = "off";
defparam \src_data[109] .lut_mask = 64'h0537053705370537;
defparam \src_data[109] .shared_arith = "off";

cyclonev_lcell_comb \src_data[110] (
	.dataa(!h2f_ARID_5),
	.datab(!h2f_AWID_5),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_110),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[110] .extended_lut = "off";
defparam \src_data[110] .lut_mask = 64'h0537053705370537;
defparam \src_data[110] .shared_arith = "off";

cyclonev_lcell_comb \src_data[111] (
	.dataa(!h2f_ARID_6),
	.datab(!h2f_AWID_6),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_111),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[111] .extended_lut = "off";
defparam \src_data[111] .lut_mask = 64'h0537053705370537;
defparam \src_data[111] .shared_arith = "off";

cyclonev_lcell_comb \src_data[112] (
	.dataa(!h2f_ARID_7),
	.datab(!h2f_AWID_7),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_112),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[112] .extended_lut = "off";
defparam \src_data[112] .lut_mask = 64'h0537053705370537;
defparam \src_data[112] .shared_arith = "off";

cyclonev_lcell_comb \src_data[113] (
	.dataa(!h2f_ARID_8),
	.datab(!h2f_AWID_8),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_113),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[113] .extended_lut = "off";
defparam \src_data[113] .lut_mask = 64'h0537053705370537;
defparam \src_data[113] .shared_arith = "off";

cyclonev_lcell_comb \src_data[114] (
	.dataa(!h2f_ARID_9),
	.datab(!h2f_AWID_9),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_114),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[114] .extended_lut = "off";
defparam \src_data[114] .lut_mask = 64'h0537053705370537;
defparam \src_data[114] .shared_arith = "off";

cyclonev_lcell_comb \src_data[115] (
	.dataa(!h2f_ARID_10),
	.datab(!h2f_AWID_10),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_115),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[115] .extended_lut = "off";
defparam \src_data[115] .lut_mask = 64'h0537053705370537;
defparam \src_data[115] .shared_arith = "off";

cyclonev_lcell_comb \src_data[116] (
	.dataa(!h2f_ARID_11),
	.datab(!h2f_AWID_11),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_116),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[116] .extended_lut = "off";
defparam \src_data[116] .lut_mask = 64'h0537053705370537;
defparam \src_data[116] .shared_arith = "off";

cyclonev_lcell_comb \src_data[86] (
	.dataa(!h2f_ARSIZE_0),
	.datab(!h2f_AWSIZE_0),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_86),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[86] .extended_lut = "off";
defparam \src_data[86] .lut_mask = 64'h0537053705370537;
defparam \src_data[86] .shared_arith = "off";

cyclonev_lcell_comb \src_data[80] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector5),
	.datad(!Selector12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_80),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[80] .extended_lut = "off";
defparam \src_data[80] .lut_mask = 64'h0357035703570357;
defparam \src_data[80] .shared_arith = "off";

cyclonev_lcell_comb \src_data[79] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector6),
	.datad(!Selector13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_79),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[79] .extended_lut = "off";
defparam \src_data[79] .lut_mask = 64'h0357035703570357;
defparam \src_data[79] .shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!\update_grant~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \update_grant~0 (
	.dataa(!nxt_in_ready1),
	.datab(!nxt_in_ready),
	.datac(!src_valid),
	.datad(!src_valid1),
	.datae(!src_payload_0),
	.dataf(!\packet_in_progress~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\update_grant~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \update_grant~0 .extended_lut = "off";
defparam \update_grant~0 .lut_mask = 64'hF000F77700000777;
defparam \update_grant~0 .shared_arith = "off";

cyclonev_lcell_comb \src_valid~0 (
	.dataa(!h2f_ARVALID_0),
	.datab(!h2f_ARADDR_4),
	.datac(!h2f_ARADDR_5),
	.datad(!h2f_ARADDR_6),
	.datae(!h2f_ARADDR_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~0 .extended_lut = "off";
defparam \src_valid~0 .lut_mask = 64'h0010000000100000;
defparam \src_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src_valid~1 (
	.dataa(!h2f_ARADDR_7),
	.datab(!has_pending_responses),
	.datac(!last_channel_13),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_valid~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~1 .extended_lut = "off";
defparam \src_valid~1 .lut_mask = 64'h4545454545454545;
defparam \src_valid~1 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_arbitrator_12 (
	nxt_in_ready,
	nxt_in_ready1,
	Equal13,
	reset,
	Equal5,
	src13_valid,
	src_payload_0,
	src13_valid1,
	src_valid,
	grant_1,
	packet_in_progress,
	grant_0,
	WideOr1,
	clk)/* synthesis synthesis_greybox=0 */;
input 	nxt_in_ready;
input 	nxt_in_ready1;
input 	Equal13;
input 	reset;
input 	Equal5;
input 	src13_valid;
input 	src_payload_0;
input 	src13_valid1;
input 	src_valid;
output 	grant_1;
input 	packet_in_progress;
output 	grant_0;
input 	WideOr1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg[0]~2_combout ;
wire \top_priority_reg[0]~q ;


cyclonev_lcell_comb \grant[1]~0 (
	.dataa(!\top_priority_reg[1]~q ),
	.datab(!\top_priority_reg[0]~q ),
	.datac(!src13_valid1),
	.datad(!src_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[1]~0 .extended_lut = "off";
defparam \grant[1]~0 .lut_mask = 64'h00D500D500D500D5;
defparam \grant[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \grant[0]~1 (
	.dataa(!\top_priority_reg[1]~q ),
	.datab(!\top_priority_reg[0]~q ),
	.datac(!src13_valid1),
	.datad(!src_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[0]~1 .extended_lut = "off";
defparam \grant[0]~1 .lut_mask = 64'h0D0C0D0C0D0C0D0C;
defparam \grant[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~0 (
	.dataa(!Equal5),
	.datab(!Equal13),
	.datac(!src13_valid),
	.datad(!src_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~0 .extended_lut = "off";
defparam \top_priority_reg[0]~0 .lut_mask = 64'hFE00FE00FE00FE00;
defparam \top_priority_reg[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~1 (
	.dataa(!nxt_in_ready1),
	.datab(!nxt_in_ready),
	.datac(!WideOr1),
	.datad(!src_payload_0),
	.datae(!packet_in_progress),
	.dataf(!\top_priority_reg[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~1 .extended_lut = "off";
defparam \top_priority_reg[0]~1 .lut_mask = 64'h0F7F007000000000;
defparam \top_priority_reg[0]~1 .shared_arith = "off";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~1_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

cyclonev_lcell_comb \top_priority_reg[0]~2 (
	.dataa(!grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~2 .extended_lut = "off";
defparam \top_priority_reg[0]~2 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \top_priority_reg[0]~2 .shared_arith = "off";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~1_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

endmodule

module spw_babasu_spw_babasu_mm_interconnect_0_cmd_mux_14 (
	h2f_WLAST_0,
	h2f_ARID_0,
	h2f_ARID_1,
	h2f_ARID_2,
	h2f_ARID_3,
	h2f_ARID_4,
	h2f_ARID_5,
	h2f_ARID_6,
	h2f_ARID_7,
	h2f_ARID_8,
	h2f_ARID_9,
	h2f_ARID_10,
	h2f_ARID_11,
	h2f_ARSIZE_0,
	h2f_ARSIZE_1,
	h2f_ARSIZE_2,
	h2f_AWID_0,
	h2f_AWID_1,
	h2f_AWID_2,
	h2f_AWID_3,
	h2f_AWID_4,
	h2f_AWID_5,
	h2f_AWID_6,
	h2f_AWID_7,
	h2f_AWID_8,
	h2f_AWID_9,
	h2f_AWID_10,
	h2f_AWID_11,
	h2f_AWSIZE_0,
	h2f_AWSIZE_1,
	h2f_AWSIZE_2,
	h2f_WDATA_0,
	h2f_WDATA_1,
	h2f_WDATA_2,
	h2f_WDATA_3,
	h2f_WDATA_4,
	h2f_WDATA_5,
	h2f_WDATA_6,
	h2f_WDATA_7,
	h2f_WSTRB_0,
	h2f_WSTRB_1,
	h2f_WSTRB_2,
	h2f_WSTRB_3,
	nxt_in_ready,
	nxt_in_ready1,
	saved_grant_1,
	Equal14,
	write_addr_data_both_valid,
	out_data_4,
	Equal141,
	Equal13,
	saved_grant_0,
	altera_reset_synchronizer_int_chain_out,
	Equal142,
	src14_valid,
	src14_valid1,
	src14_valid2,
	src_valid,
	src_data_87,
	src_data_88,
	src_valid1,
	src_data_35,
	src_data_34,
	src_data_33,
	src_data_32,
	src_payload_0,
	src14_valid3,
	src14_valid4,
	Selector3,
	Selector10,
	Selector4,
	Selector11,
	src_payload,
	src_data_82,
	src_data_81,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_data_105,
	src_data_106,
	src_data_107,
	src_data_108,
	src_data_109,
	src_data_110,
	src_data_111,
	src_data_112,
	src_data_113,
	src_data_114,
	src_data_115,
	src_data_116,
	src_data_86,
	Selector5,
	Selector12,
	src_data_80,
	Selector6,
	Selector13,
	src_data_79,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_WLAST_0;
input 	h2f_ARID_0;
input 	h2f_ARID_1;
input 	h2f_ARID_2;
input 	h2f_ARID_3;
input 	h2f_ARID_4;
input 	h2f_ARID_5;
input 	h2f_ARID_6;
input 	h2f_ARID_7;
input 	h2f_ARID_8;
input 	h2f_ARID_9;
input 	h2f_ARID_10;
input 	h2f_ARID_11;
input 	h2f_ARSIZE_0;
input 	h2f_ARSIZE_1;
input 	h2f_ARSIZE_2;
input 	h2f_AWID_0;
input 	h2f_AWID_1;
input 	h2f_AWID_2;
input 	h2f_AWID_3;
input 	h2f_AWID_4;
input 	h2f_AWID_5;
input 	h2f_AWID_6;
input 	h2f_AWID_7;
input 	h2f_AWID_8;
input 	h2f_AWID_9;
input 	h2f_AWID_10;
input 	h2f_AWID_11;
input 	h2f_AWSIZE_0;
input 	h2f_AWSIZE_1;
input 	h2f_AWSIZE_2;
input 	h2f_WDATA_0;
input 	h2f_WDATA_1;
input 	h2f_WDATA_2;
input 	h2f_WDATA_3;
input 	h2f_WDATA_4;
input 	h2f_WDATA_5;
input 	h2f_WDATA_6;
input 	h2f_WDATA_7;
input 	h2f_WSTRB_0;
input 	h2f_WSTRB_1;
input 	h2f_WSTRB_2;
input 	h2f_WSTRB_3;
input 	nxt_in_ready;
input 	nxt_in_ready1;
output 	saved_grant_1;
input 	Equal14;
input 	write_addr_data_both_valid;
input 	out_data_4;
input 	Equal141;
input 	Equal13;
output 	saved_grant_0;
input 	altera_reset_synchronizer_int_chain_out;
input 	Equal142;
input 	src14_valid;
input 	src14_valid1;
input 	src14_valid2;
output 	src_valid;
output 	src_data_87;
output 	src_data_88;
output 	src_valid1;
output 	src_data_35;
output 	src_data_34;
output 	src_data_33;
output 	src_data_32;
output 	src_payload_0;
input 	src14_valid3;
input 	src14_valid4;
input 	Selector3;
input 	Selector10;
input 	Selector4;
input 	Selector11;
output 	src_payload;
output 	src_data_82;
output 	src_data_81;
output 	src_payload1;
output 	src_payload2;
output 	src_payload3;
output 	src_payload4;
output 	src_payload5;
output 	src_payload6;
output 	src_payload7;
output 	src_data_105;
output 	src_data_106;
output 	src_data_107;
output 	src_data_108;
output 	src_data_109;
output 	src_data_110;
output 	src_data_111;
output 	src_data_112;
output 	src_data_113;
output 	src_data_114;
output 	src_data_115;
output 	src_data_116;
output 	src_data_86;
input 	Selector5;
input 	Selector12;
output 	src_data_80;
input 	Selector6;
input 	Selector13;
output 	src_data_79;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[1]~0_combout ;
wire \arb|grant[0]~1_combout ;
wire \WideOr1~combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~0_combout ;


spw_babasu_altera_merlin_arbitrator_13 arb(
	.nxt_in_ready(nxt_in_ready),
	.nxt_in_ready1(nxt_in_ready1),
	.Equal13(Equal13),
	.reset(altera_reset_synchronizer_int_chain_out),
	.Equal14(Equal142),
	.src14_valid(src14_valid1),
	.src_payload_0(src_payload_0),
	.src14_valid1(src14_valid3),
	.src14_valid2(src14_valid4),
	.grant_1(\arb|grant[1]~0_combout ),
	.packet_in_progress(\packet_in_progress~q ),
	.grant_0(\arb|grant[0]~1_combout ),
	.WideOr1(\WideOr1~combout ),
	.clk(clk_clk));

cyclonev_lcell_comb WideOr1(
	.dataa(!Equal142),
	.datab(!Equal13),
	.datac(!saved_grant_0),
	.datad(!src14_valid1),
	.datae(!src_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr1.extended_lut = "off";
defparam WideOr1.lut_mask = 64'hFFFE0000FFFE0000;
defparam WideOr1.shared_arith = "off";

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

cyclonev_lcell_comb \src_valid~0 (
	.dataa(!saved_grant_1),
	.datab(!Equal14),
	.datac(!src14_valid2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~0 .extended_lut = "off";
defparam \src_valid~0 .lut_mask = 64'h0101010101010101;
defparam \src_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[87] (
	.dataa(!h2f_ARSIZE_1),
	.datab(!h2f_AWSIZE_1),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_87),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[87] .extended_lut = "off";
defparam \src_data[87] .lut_mask = 64'h0537053705370537;
defparam \src_data[87] .shared_arith = "off";

cyclonev_lcell_comb \src_data[88] (
	.dataa(!h2f_ARSIZE_2),
	.datab(!h2f_AWSIZE_2),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_88),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[88] .extended_lut = "off";
defparam \src_data[88] .lut_mask = 64'h0537053705370537;
defparam \src_data[88] .shared_arith = "off";

cyclonev_lcell_comb \src_valid~1 (
	.dataa(!out_data_4),
	.datab(!Equal141),
	.datac(!Equal13),
	.datad(!saved_grant_0),
	.datae(!write_addr_data_both_valid),
	.dataf(!src14_valid),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~1 .extended_lut = "off";
defparam \src_valid~1 .lut_mask = 64'h0000000200000000;
defparam \src_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \src_data[35] (
	.dataa(!h2f_WSTRB_3),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_35),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[35] .extended_lut = "off";
defparam \src_data[35] .lut_mask = 64'h3737373737373737;
defparam \src_data[35] .shared_arith = "off";

cyclonev_lcell_comb \src_data[34] (
	.dataa(!h2f_WSTRB_2),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_34),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[34] .extended_lut = "off";
defparam \src_data[34] .lut_mask = 64'h3737373737373737;
defparam \src_data[34] .shared_arith = "off";

cyclonev_lcell_comb \src_data[33] (
	.dataa(!h2f_WSTRB_1),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_33),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[33] .extended_lut = "off";
defparam \src_data[33] .lut_mask = 64'h3737373737373737;
defparam \src_data[33] .shared_arith = "off";

cyclonev_lcell_comb \src_data[32] (
	.dataa(!h2f_WSTRB_0),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_32),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[32] .extended_lut = "off";
defparam \src_data[32] .lut_mask = 64'h3737373737373737;
defparam \src_data[32] .shared_arith = "off";

cyclonev_lcell_comb \src_payload[0] (
	.dataa(!h2f_WLAST_0),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload[0] .extended_lut = "off";
defparam \src_payload[0] .lut_mask = 64'h3737373737373737;
defparam \src_payload[0] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!h2f_WDATA_0),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h1111111111111111;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[82] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector3),
	.datad(!Selector10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_82),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[82] .extended_lut = "off";
defparam \src_data[82] .lut_mask = 64'h0357035703570357;
defparam \src_data[82] .shared_arith = "off";

cyclonev_lcell_comb \src_data[81] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector4),
	.datad(!Selector11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_81),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[81] .extended_lut = "off";
defparam \src_data[81] .lut_mask = 64'h0357035703570357;
defparam \src_data[81] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!h2f_WDATA_1),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h1111111111111111;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!h2f_WDATA_2),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h1111111111111111;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~3 (
	.dataa(!h2f_WDATA_3),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~3 .extended_lut = "off";
defparam \src_payload~3 .lut_mask = 64'h1111111111111111;
defparam \src_payload~3 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~4 (
	.dataa(!h2f_WDATA_4),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~4 .extended_lut = "off";
defparam \src_payload~4 .lut_mask = 64'h1111111111111111;
defparam \src_payload~4 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~5 (
	.dataa(!h2f_WDATA_5),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~5 .extended_lut = "off";
defparam \src_payload~5 .lut_mask = 64'h1111111111111111;
defparam \src_payload~5 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~6 (
	.dataa(!h2f_WDATA_6),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~6 .extended_lut = "off";
defparam \src_payload~6 .lut_mask = 64'h1111111111111111;
defparam \src_payload~6 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~7 (
	.dataa(!h2f_WDATA_7),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~7 .extended_lut = "off";
defparam \src_payload~7 .lut_mask = 64'h1111111111111111;
defparam \src_payload~7 .shared_arith = "off";

cyclonev_lcell_comb \src_data[105] (
	.dataa(!h2f_ARID_0),
	.datab(!h2f_AWID_0),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_105),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[105] .extended_lut = "off";
defparam \src_data[105] .lut_mask = 64'h0537053705370537;
defparam \src_data[105] .shared_arith = "off";

cyclonev_lcell_comb \src_data[106] (
	.dataa(!h2f_ARID_1),
	.datab(!h2f_AWID_1),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_106),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[106] .extended_lut = "off";
defparam \src_data[106] .lut_mask = 64'h0537053705370537;
defparam \src_data[106] .shared_arith = "off";

cyclonev_lcell_comb \src_data[107] (
	.dataa(!h2f_ARID_2),
	.datab(!h2f_AWID_2),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_107),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[107] .extended_lut = "off";
defparam \src_data[107] .lut_mask = 64'h0537053705370537;
defparam \src_data[107] .shared_arith = "off";

cyclonev_lcell_comb \src_data[108] (
	.dataa(!h2f_ARID_3),
	.datab(!h2f_AWID_3),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_108),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[108] .extended_lut = "off";
defparam \src_data[108] .lut_mask = 64'h0537053705370537;
defparam \src_data[108] .shared_arith = "off";

cyclonev_lcell_comb \src_data[109] (
	.dataa(!h2f_ARID_4),
	.datab(!h2f_AWID_4),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_109),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[109] .extended_lut = "off";
defparam \src_data[109] .lut_mask = 64'h0537053705370537;
defparam \src_data[109] .shared_arith = "off";

cyclonev_lcell_comb \src_data[110] (
	.dataa(!h2f_ARID_5),
	.datab(!h2f_AWID_5),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_110),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[110] .extended_lut = "off";
defparam \src_data[110] .lut_mask = 64'h0537053705370537;
defparam \src_data[110] .shared_arith = "off";

cyclonev_lcell_comb \src_data[111] (
	.dataa(!h2f_ARID_6),
	.datab(!h2f_AWID_6),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_111),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[111] .extended_lut = "off";
defparam \src_data[111] .lut_mask = 64'h0537053705370537;
defparam \src_data[111] .shared_arith = "off";

cyclonev_lcell_comb \src_data[112] (
	.dataa(!h2f_ARID_7),
	.datab(!h2f_AWID_7),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_112),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[112] .extended_lut = "off";
defparam \src_data[112] .lut_mask = 64'h0537053705370537;
defparam \src_data[112] .shared_arith = "off";

cyclonev_lcell_comb \src_data[113] (
	.dataa(!h2f_ARID_8),
	.datab(!h2f_AWID_8),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_113),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[113] .extended_lut = "off";
defparam \src_data[113] .lut_mask = 64'h0537053705370537;
defparam \src_data[113] .shared_arith = "off";

cyclonev_lcell_comb \src_data[114] (
	.dataa(!h2f_ARID_9),
	.datab(!h2f_AWID_9),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_114),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[114] .extended_lut = "off";
defparam \src_data[114] .lut_mask = 64'h0537053705370537;
defparam \src_data[114] .shared_arith = "off";

cyclonev_lcell_comb \src_data[115] (
	.dataa(!h2f_ARID_10),
	.datab(!h2f_AWID_10),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_115),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[115] .extended_lut = "off";
defparam \src_data[115] .lut_mask = 64'h0537053705370537;
defparam \src_data[115] .shared_arith = "off";

cyclonev_lcell_comb \src_data[116] (
	.dataa(!h2f_ARID_11),
	.datab(!h2f_AWID_11),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_116),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[116] .extended_lut = "off";
defparam \src_data[116] .lut_mask = 64'h0537053705370537;
defparam \src_data[116] .shared_arith = "off";

cyclonev_lcell_comb \src_data[86] (
	.dataa(!h2f_ARSIZE_0),
	.datab(!h2f_AWSIZE_0),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_86),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[86] .extended_lut = "off";
defparam \src_data[86] .lut_mask = 64'h0537053705370537;
defparam \src_data[86] .shared_arith = "off";

cyclonev_lcell_comb \src_data[80] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector5),
	.datad(!Selector12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_80),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[80] .extended_lut = "off";
defparam \src_data[80] .lut_mask = 64'h0357035703570357;
defparam \src_data[80] .shared_arith = "off";

cyclonev_lcell_comb \src_data[79] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector6),
	.datad(!Selector13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_79),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[79] .extended_lut = "off";
defparam \src_data[79] .lut_mask = 64'h0357035703570357;
defparam \src_data[79] .shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!\update_grant~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \update_grant~0 (
	.dataa(!nxt_in_ready1),
	.datab(!nxt_in_ready),
	.datac(!src_valid),
	.datad(!src_valid1),
	.datae(!src_payload_0),
	.dataf(!\packet_in_progress~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\update_grant~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \update_grant~0 .extended_lut = "off";
defparam \update_grant~0 .lut_mask = 64'hF000F77700000777;
defparam \update_grant~0 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_arbitrator_13 (
	nxt_in_ready,
	nxt_in_ready1,
	Equal13,
	reset,
	Equal14,
	src14_valid,
	src_payload_0,
	src14_valid1,
	src14_valid2,
	grant_1,
	packet_in_progress,
	grant_0,
	WideOr1,
	clk)/* synthesis synthesis_greybox=0 */;
input 	nxt_in_ready;
input 	nxt_in_ready1;
input 	Equal13;
input 	reset;
input 	Equal14;
input 	src14_valid;
input 	src_payload_0;
input 	src14_valid1;
input 	src14_valid2;
output 	grant_1;
input 	packet_in_progress;
output 	grant_0;
input 	WideOr1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg[0]~2_combout ;
wire \top_priority_reg[0]~q ;


cyclonev_lcell_comb \grant[1]~0 (
	.dataa(!\top_priority_reg[1]~q ),
	.datab(!\top_priority_reg[0]~q ),
	.datac(!src14_valid1),
	.datad(!src14_valid2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[1]~0 .extended_lut = "off";
defparam \grant[1]~0 .lut_mask = 64'h00D500D500D500D5;
defparam \grant[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \grant[0]~1 (
	.dataa(!\top_priority_reg[1]~q ),
	.datab(!\top_priority_reg[0]~q ),
	.datac(!src14_valid1),
	.datad(!src14_valid2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[0]~1 .extended_lut = "off";
defparam \grant[0]~1 .lut_mask = 64'h0D0C0D0C0D0C0D0C;
defparam \grant[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~0 (
	.dataa(!Equal14),
	.datab(!Equal13),
	.datac(!src14_valid),
	.datad(!src14_valid2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~0 .extended_lut = "off";
defparam \top_priority_reg[0]~0 .lut_mask = 64'hFE00FE00FE00FE00;
defparam \top_priority_reg[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~1 (
	.dataa(!nxt_in_ready1),
	.datab(!nxt_in_ready),
	.datac(!WideOr1),
	.datad(!src_payload_0),
	.datae(!packet_in_progress),
	.dataf(!\top_priority_reg[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~1 .extended_lut = "off";
defparam \top_priority_reg[0]~1 .lut_mask = 64'h0F7F007000000000;
defparam \top_priority_reg[0]~1 .shared_arith = "off";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~1_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

cyclonev_lcell_comb \top_priority_reg[0]~2 (
	.dataa(!grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~2 .extended_lut = "off";
defparam \top_priority_reg[0]~2 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \top_priority_reg[0]~2 .shared_arith = "off";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~1_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

endmodule

module spw_babasu_spw_babasu_mm_interconnect_0_cmd_mux_15 (
	h2f_WLAST_0,
	h2f_ARID_0,
	h2f_ARID_1,
	h2f_ARID_2,
	h2f_ARID_3,
	h2f_ARID_4,
	h2f_ARID_5,
	h2f_ARID_6,
	h2f_ARID_7,
	h2f_ARID_8,
	h2f_ARID_9,
	h2f_ARID_10,
	h2f_ARID_11,
	h2f_ARSIZE_0,
	h2f_ARSIZE_1,
	h2f_ARSIZE_2,
	h2f_AWID_0,
	h2f_AWID_1,
	h2f_AWID_2,
	h2f_AWID_3,
	h2f_AWID_4,
	h2f_AWID_5,
	h2f_AWID_6,
	h2f_AWID_7,
	h2f_AWID_8,
	h2f_AWID_9,
	h2f_AWID_10,
	h2f_AWID_11,
	h2f_AWSIZE_0,
	h2f_AWSIZE_1,
	h2f_AWSIZE_2,
	h2f_WDATA_0,
	h2f_WDATA_1,
	h2f_WDATA_2,
	h2f_WDATA_3,
	h2f_WDATA_4,
	h2f_WDATA_5,
	h2f_WDATA_6,
	h2f_WSTRB_0,
	h2f_WSTRB_1,
	h2f_WSTRB_2,
	h2f_WSTRB_3,
	nxt_in_ready,
	nxt_in_ready1,
	saved_grant_1,
	Equal15,
	write_addr_data_both_valid,
	out_data_5,
	Equal13,
	Equal151,
	saved_grant_0,
	altera_reset_synchronizer_int_chain_out,
	Equal152,
	src15_valid,
	src15_valid1,
	src15_valid2,
	src_valid,
	src_data_87,
	src_data_88,
	src_valid1,
	src_data_35,
	src_data_34,
	src_data_33,
	src_data_32,
	src_payload_0,
	src15_valid3,
	src15_valid4,
	Selector3,
	Selector10,
	Selector4,
	Selector11,
	src_payload,
	src_data_82,
	src_data_81,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_data_105,
	src_data_106,
	src_data_107,
	src_data_108,
	src_data_109,
	src_data_110,
	src_data_111,
	src_data_112,
	src_data_113,
	src_data_114,
	src_data_115,
	src_data_116,
	src_data_86,
	Selector5,
	Selector12,
	src_data_80,
	Selector6,
	Selector13,
	src_data_79,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_WLAST_0;
input 	h2f_ARID_0;
input 	h2f_ARID_1;
input 	h2f_ARID_2;
input 	h2f_ARID_3;
input 	h2f_ARID_4;
input 	h2f_ARID_5;
input 	h2f_ARID_6;
input 	h2f_ARID_7;
input 	h2f_ARID_8;
input 	h2f_ARID_9;
input 	h2f_ARID_10;
input 	h2f_ARID_11;
input 	h2f_ARSIZE_0;
input 	h2f_ARSIZE_1;
input 	h2f_ARSIZE_2;
input 	h2f_AWID_0;
input 	h2f_AWID_1;
input 	h2f_AWID_2;
input 	h2f_AWID_3;
input 	h2f_AWID_4;
input 	h2f_AWID_5;
input 	h2f_AWID_6;
input 	h2f_AWID_7;
input 	h2f_AWID_8;
input 	h2f_AWID_9;
input 	h2f_AWID_10;
input 	h2f_AWID_11;
input 	h2f_AWSIZE_0;
input 	h2f_AWSIZE_1;
input 	h2f_AWSIZE_2;
input 	h2f_WDATA_0;
input 	h2f_WDATA_1;
input 	h2f_WDATA_2;
input 	h2f_WDATA_3;
input 	h2f_WDATA_4;
input 	h2f_WDATA_5;
input 	h2f_WDATA_6;
input 	h2f_WSTRB_0;
input 	h2f_WSTRB_1;
input 	h2f_WSTRB_2;
input 	h2f_WSTRB_3;
input 	nxt_in_ready;
input 	nxt_in_ready1;
output 	saved_grant_1;
input 	Equal15;
input 	write_addr_data_both_valid;
input 	out_data_5;
input 	Equal13;
input 	Equal151;
output 	saved_grant_0;
input 	altera_reset_synchronizer_int_chain_out;
input 	Equal152;
input 	src15_valid;
input 	src15_valid1;
input 	src15_valid2;
output 	src_valid;
output 	src_data_87;
output 	src_data_88;
output 	src_valid1;
output 	src_data_35;
output 	src_data_34;
output 	src_data_33;
output 	src_data_32;
output 	src_payload_0;
input 	src15_valid3;
input 	src15_valid4;
input 	Selector3;
input 	Selector10;
input 	Selector4;
input 	Selector11;
output 	src_payload;
output 	src_data_82;
output 	src_data_81;
output 	src_payload1;
output 	src_payload2;
output 	src_payload3;
output 	src_payload4;
output 	src_payload5;
output 	src_payload6;
output 	src_data_105;
output 	src_data_106;
output 	src_data_107;
output 	src_data_108;
output 	src_data_109;
output 	src_data_110;
output 	src_data_111;
output 	src_data_112;
output 	src_data_113;
output 	src_data_114;
output 	src_data_115;
output 	src_data_116;
output 	src_data_86;
input 	Selector5;
input 	Selector12;
output 	src_data_80;
input 	Selector6;
input 	Selector13;
output 	src_data_79;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[1]~0_combout ;
wire \arb|grant[0]~1_combout ;
wire \WideOr1~combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~0_combout ;


spw_babasu_altera_merlin_arbitrator_14 arb(
	.nxt_in_ready(nxt_in_ready),
	.nxt_in_ready1(nxt_in_ready1),
	.Equal15(Equal151),
	.reset(altera_reset_synchronizer_int_chain_out),
	.Equal151(Equal152),
	.src15_valid(src15_valid1),
	.src_payload_0(src_payload_0),
	.src15_valid1(src15_valid3),
	.src15_valid2(src15_valid4),
	.grant_1(\arb|grant[1]~0_combout ),
	.packet_in_progress(\packet_in_progress~q ),
	.grant_0(\arb|grant[0]~1_combout ),
	.WideOr1(\WideOr1~combout ),
	.clk(clk_clk));

cyclonev_lcell_comb WideOr1(
	.dataa(!Equal151),
	.datab(!Equal152),
	.datac(!saved_grant_0),
	.datad(!src15_valid1),
	.datae(!src_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr1.extended_lut = "off";
defparam WideOr1.lut_mask = 64'hFFFE0000FFFE0000;
defparam WideOr1.shared_arith = "off";

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

cyclonev_lcell_comb \src_valid~0 (
	.dataa(!saved_grant_1),
	.datab(!Equal15),
	.datac(!src15_valid2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~0 .extended_lut = "off";
defparam \src_valid~0 .lut_mask = 64'h0101010101010101;
defparam \src_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[87] (
	.dataa(!h2f_ARSIZE_1),
	.datab(!h2f_AWSIZE_1),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_87),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[87] .extended_lut = "off";
defparam \src_data[87] .lut_mask = 64'h0537053705370537;
defparam \src_data[87] .shared_arith = "off";

cyclonev_lcell_comb \src_data[88] (
	.dataa(!h2f_ARSIZE_2),
	.datab(!h2f_AWSIZE_2),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_88),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[88] .extended_lut = "off";
defparam \src_data[88] .lut_mask = 64'h0537053705370537;
defparam \src_data[88] .shared_arith = "off";

cyclonev_lcell_comb \src_valid~1 (
	.dataa(!out_data_5),
	.datab(!Equal151),
	.datac(!Equal13),
	.datad(!saved_grant_0),
	.datae(!write_addr_data_both_valid),
	.dataf(!src15_valid),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~1 .extended_lut = "off";
defparam \src_valid~1 .lut_mask = 64'h0000000100000000;
defparam \src_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \src_data[35] (
	.dataa(!h2f_WSTRB_3),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_35),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[35] .extended_lut = "off";
defparam \src_data[35] .lut_mask = 64'h3737373737373737;
defparam \src_data[35] .shared_arith = "off";

cyclonev_lcell_comb \src_data[34] (
	.dataa(!h2f_WSTRB_2),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_34),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[34] .extended_lut = "off";
defparam \src_data[34] .lut_mask = 64'h3737373737373737;
defparam \src_data[34] .shared_arith = "off";

cyclonev_lcell_comb \src_data[33] (
	.dataa(!h2f_WSTRB_1),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_33),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[33] .extended_lut = "off";
defparam \src_data[33] .lut_mask = 64'h3737373737373737;
defparam \src_data[33] .shared_arith = "off";

cyclonev_lcell_comb \src_data[32] (
	.dataa(!h2f_WSTRB_0),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_32),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[32] .extended_lut = "off";
defparam \src_data[32] .lut_mask = 64'h3737373737373737;
defparam \src_data[32] .shared_arith = "off";

cyclonev_lcell_comb \src_payload[0] (
	.dataa(!h2f_WLAST_0),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload[0] .extended_lut = "off";
defparam \src_payload[0] .lut_mask = 64'h3737373737373737;
defparam \src_payload[0] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!h2f_WDATA_0),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h1111111111111111;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[82] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector3),
	.datad(!Selector10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_82),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[82] .extended_lut = "off";
defparam \src_data[82] .lut_mask = 64'h0357035703570357;
defparam \src_data[82] .shared_arith = "off";

cyclonev_lcell_comb \src_data[81] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector4),
	.datad(!Selector11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_81),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[81] .extended_lut = "off";
defparam \src_data[81] .lut_mask = 64'h0357035703570357;
defparam \src_data[81] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!h2f_WDATA_1),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h1111111111111111;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!h2f_WDATA_2),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h1111111111111111;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~3 (
	.dataa(!h2f_WDATA_3),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~3 .extended_lut = "off";
defparam \src_payload~3 .lut_mask = 64'h1111111111111111;
defparam \src_payload~3 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~4 (
	.dataa(!h2f_WDATA_4),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~4 .extended_lut = "off";
defparam \src_payload~4 .lut_mask = 64'h1111111111111111;
defparam \src_payload~4 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~5 (
	.dataa(!h2f_WDATA_5),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~5 .extended_lut = "off";
defparam \src_payload~5 .lut_mask = 64'h1111111111111111;
defparam \src_payload~5 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~6 (
	.dataa(!h2f_WDATA_6),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~6 .extended_lut = "off";
defparam \src_payload~6 .lut_mask = 64'h1111111111111111;
defparam \src_payload~6 .shared_arith = "off";

cyclonev_lcell_comb \src_data[105] (
	.dataa(!h2f_ARID_0),
	.datab(!h2f_AWID_0),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_105),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[105] .extended_lut = "off";
defparam \src_data[105] .lut_mask = 64'h0537053705370537;
defparam \src_data[105] .shared_arith = "off";

cyclonev_lcell_comb \src_data[106] (
	.dataa(!h2f_ARID_1),
	.datab(!h2f_AWID_1),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_106),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[106] .extended_lut = "off";
defparam \src_data[106] .lut_mask = 64'h0537053705370537;
defparam \src_data[106] .shared_arith = "off";

cyclonev_lcell_comb \src_data[107] (
	.dataa(!h2f_ARID_2),
	.datab(!h2f_AWID_2),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_107),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[107] .extended_lut = "off";
defparam \src_data[107] .lut_mask = 64'h0537053705370537;
defparam \src_data[107] .shared_arith = "off";

cyclonev_lcell_comb \src_data[108] (
	.dataa(!h2f_ARID_3),
	.datab(!h2f_AWID_3),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_108),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[108] .extended_lut = "off";
defparam \src_data[108] .lut_mask = 64'h0537053705370537;
defparam \src_data[108] .shared_arith = "off";

cyclonev_lcell_comb \src_data[109] (
	.dataa(!h2f_ARID_4),
	.datab(!h2f_AWID_4),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_109),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[109] .extended_lut = "off";
defparam \src_data[109] .lut_mask = 64'h0537053705370537;
defparam \src_data[109] .shared_arith = "off";

cyclonev_lcell_comb \src_data[110] (
	.dataa(!h2f_ARID_5),
	.datab(!h2f_AWID_5),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_110),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[110] .extended_lut = "off";
defparam \src_data[110] .lut_mask = 64'h0537053705370537;
defparam \src_data[110] .shared_arith = "off";

cyclonev_lcell_comb \src_data[111] (
	.dataa(!h2f_ARID_6),
	.datab(!h2f_AWID_6),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_111),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[111] .extended_lut = "off";
defparam \src_data[111] .lut_mask = 64'h0537053705370537;
defparam \src_data[111] .shared_arith = "off";

cyclonev_lcell_comb \src_data[112] (
	.dataa(!h2f_ARID_7),
	.datab(!h2f_AWID_7),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_112),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[112] .extended_lut = "off";
defparam \src_data[112] .lut_mask = 64'h0537053705370537;
defparam \src_data[112] .shared_arith = "off";

cyclonev_lcell_comb \src_data[113] (
	.dataa(!h2f_ARID_8),
	.datab(!h2f_AWID_8),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_113),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[113] .extended_lut = "off";
defparam \src_data[113] .lut_mask = 64'h0537053705370537;
defparam \src_data[113] .shared_arith = "off";

cyclonev_lcell_comb \src_data[114] (
	.dataa(!h2f_ARID_9),
	.datab(!h2f_AWID_9),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_114),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[114] .extended_lut = "off";
defparam \src_data[114] .lut_mask = 64'h0537053705370537;
defparam \src_data[114] .shared_arith = "off";

cyclonev_lcell_comb \src_data[115] (
	.dataa(!h2f_ARID_10),
	.datab(!h2f_AWID_10),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_115),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[115] .extended_lut = "off";
defparam \src_data[115] .lut_mask = 64'h0537053705370537;
defparam \src_data[115] .shared_arith = "off";

cyclonev_lcell_comb \src_data[116] (
	.dataa(!h2f_ARID_11),
	.datab(!h2f_AWID_11),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_116),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[116] .extended_lut = "off";
defparam \src_data[116] .lut_mask = 64'h0537053705370537;
defparam \src_data[116] .shared_arith = "off";

cyclonev_lcell_comb \src_data[86] (
	.dataa(!h2f_ARSIZE_0),
	.datab(!h2f_AWSIZE_0),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_86),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[86] .extended_lut = "off";
defparam \src_data[86] .lut_mask = 64'h0537053705370537;
defparam \src_data[86] .shared_arith = "off";

cyclonev_lcell_comb \src_data[80] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector5),
	.datad(!Selector12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_80),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[80] .extended_lut = "off";
defparam \src_data[80] .lut_mask = 64'h0357035703570357;
defparam \src_data[80] .shared_arith = "off";

cyclonev_lcell_comb \src_data[79] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector6),
	.datad(!Selector13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_79),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[79] .extended_lut = "off";
defparam \src_data[79] .lut_mask = 64'h0357035703570357;
defparam \src_data[79] .shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!\update_grant~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \update_grant~0 (
	.dataa(!nxt_in_ready1),
	.datab(!nxt_in_ready),
	.datac(!src_valid),
	.datad(!src_valid1),
	.datae(!src_payload_0),
	.dataf(!\packet_in_progress~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\update_grant~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \update_grant~0 .extended_lut = "off";
defparam \update_grant~0 .lut_mask = 64'hF000F77700000777;
defparam \update_grant~0 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_arbitrator_14 (
	nxt_in_ready,
	nxt_in_ready1,
	Equal15,
	reset,
	Equal151,
	src15_valid,
	src_payload_0,
	src15_valid1,
	src15_valid2,
	grant_1,
	packet_in_progress,
	grant_0,
	WideOr1,
	clk)/* synthesis synthesis_greybox=0 */;
input 	nxt_in_ready;
input 	nxt_in_ready1;
input 	Equal15;
input 	reset;
input 	Equal151;
input 	src15_valid;
input 	src_payload_0;
input 	src15_valid1;
input 	src15_valid2;
output 	grant_1;
input 	packet_in_progress;
output 	grant_0;
input 	WideOr1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg[0]~2_combout ;
wire \top_priority_reg[0]~q ;


cyclonev_lcell_comb \grant[1]~0 (
	.dataa(!\top_priority_reg[1]~q ),
	.datab(!\top_priority_reg[0]~q ),
	.datac(!src15_valid1),
	.datad(!src15_valid2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[1]~0 .extended_lut = "off";
defparam \grant[1]~0 .lut_mask = 64'h00D500D500D500D5;
defparam \grant[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \grant[0]~1 (
	.dataa(!\top_priority_reg[1]~q ),
	.datab(!\top_priority_reg[0]~q ),
	.datac(!src15_valid1),
	.datad(!src15_valid2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[0]~1 .extended_lut = "off";
defparam \grant[0]~1 .lut_mask = 64'h0D0C0D0C0D0C0D0C;
defparam \grant[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~0 (
	.dataa(!Equal15),
	.datab(!Equal151),
	.datac(!src15_valid),
	.datad(!src15_valid2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~0 .extended_lut = "off";
defparam \top_priority_reg[0]~0 .lut_mask = 64'hFE00FE00FE00FE00;
defparam \top_priority_reg[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~1 (
	.dataa(!nxt_in_ready1),
	.datab(!nxt_in_ready),
	.datac(!WideOr1),
	.datad(!src_payload_0),
	.datae(!packet_in_progress),
	.dataf(!\top_priority_reg[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~1 .extended_lut = "off";
defparam \top_priority_reg[0]~1 .lut_mask = 64'h0F7F007000000000;
defparam \top_priority_reg[0]~1 .shared_arith = "off";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~1_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

cyclonev_lcell_comb \top_priority_reg[0]~2 (
	.dataa(!grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~2 .extended_lut = "off";
defparam \top_priority_reg[0]~2 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \top_priority_reg[0]~2 .shared_arith = "off";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~1_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

endmodule

module spw_babasu_spw_babasu_mm_interconnect_0_cmd_mux_16 (
	h2f_WLAST_0,
	h2f_ARID_0,
	h2f_ARID_1,
	h2f_ARID_2,
	h2f_ARID_3,
	h2f_ARID_4,
	h2f_ARID_5,
	h2f_ARID_6,
	h2f_ARID_7,
	h2f_ARID_8,
	h2f_ARID_9,
	h2f_ARID_10,
	h2f_ARID_11,
	h2f_ARSIZE_0,
	h2f_ARSIZE_1,
	h2f_ARSIZE_2,
	h2f_AWID_0,
	h2f_AWID_1,
	h2f_AWID_2,
	h2f_AWID_3,
	h2f_AWID_4,
	h2f_AWID_5,
	h2f_AWID_6,
	h2f_AWID_7,
	h2f_AWID_8,
	h2f_AWID_9,
	h2f_AWID_10,
	h2f_AWID_11,
	h2f_AWSIZE_0,
	h2f_AWSIZE_1,
	h2f_AWSIZE_2,
	h2f_WDATA_0,
	h2f_WSTRB_0,
	h2f_WSTRB_1,
	h2f_WSTRB_2,
	h2f_WSTRB_3,
	nxt_in_ready,
	nxt_in_ready1,
	Equal16,
	saved_grant_1,
	write_addr_data_both_valid,
	out_data_4,
	Equal161,
	Equal162,
	saved_grant_0,
	altera_reset_synchronizer_int_chain_out,
	src16_valid,
	src16_valid1,
	src16_valid2,
	src_valid,
	src_valid1,
	src16_valid3,
	WideOr11,
	src_data_87,
	src_data_88,
	src_data_35,
	src_data_34,
	src_data_33,
	src_data_32,
	src_payload_0,
	src16_valid4,
	Selector3,
	Selector10,
	Selector4,
	Selector11,
	src_payload,
	src_data_82,
	src_data_81,
	src_data_105,
	src_data_106,
	src_data_107,
	src_data_108,
	src_data_109,
	src_data_110,
	src_data_111,
	src_data_112,
	src_data_113,
	src_data_114,
	src_data_115,
	src_data_116,
	src_data_86,
	Selector5,
	Selector12,
	src_data_80,
	Selector6,
	Selector13,
	src_data_79,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_WLAST_0;
input 	h2f_ARID_0;
input 	h2f_ARID_1;
input 	h2f_ARID_2;
input 	h2f_ARID_3;
input 	h2f_ARID_4;
input 	h2f_ARID_5;
input 	h2f_ARID_6;
input 	h2f_ARID_7;
input 	h2f_ARID_8;
input 	h2f_ARID_9;
input 	h2f_ARID_10;
input 	h2f_ARID_11;
input 	h2f_ARSIZE_0;
input 	h2f_ARSIZE_1;
input 	h2f_ARSIZE_2;
input 	h2f_AWID_0;
input 	h2f_AWID_1;
input 	h2f_AWID_2;
input 	h2f_AWID_3;
input 	h2f_AWID_4;
input 	h2f_AWID_5;
input 	h2f_AWID_6;
input 	h2f_AWID_7;
input 	h2f_AWID_8;
input 	h2f_AWID_9;
input 	h2f_AWID_10;
input 	h2f_AWID_11;
input 	h2f_AWSIZE_0;
input 	h2f_AWSIZE_1;
input 	h2f_AWSIZE_2;
input 	h2f_WDATA_0;
input 	h2f_WSTRB_0;
input 	h2f_WSTRB_1;
input 	h2f_WSTRB_2;
input 	h2f_WSTRB_3;
input 	nxt_in_ready;
input 	nxt_in_ready1;
input 	Equal16;
output 	saved_grant_1;
input 	write_addr_data_both_valid;
input 	out_data_4;
input 	Equal161;
input 	Equal162;
output 	saved_grant_0;
input 	altera_reset_synchronizer_int_chain_out;
input 	src16_valid;
input 	src16_valid1;
input 	src16_valid2;
output 	src_valid;
output 	src_valid1;
input 	src16_valid3;
output 	WideOr11;
output 	src_data_87;
output 	src_data_88;
output 	src_data_35;
output 	src_data_34;
output 	src_data_33;
output 	src_data_32;
output 	src_payload_0;
input 	src16_valid4;
input 	Selector3;
input 	Selector10;
input 	Selector4;
input 	Selector11;
output 	src_payload;
output 	src_data_82;
output 	src_data_81;
output 	src_data_105;
output 	src_data_106;
output 	src_data_107;
output 	src_data_108;
output 	src_data_109;
output 	src_data_110;
output 	src_data_111;
output 	src_data_112;
output 	src_data_113;
output 	src_data_114;
output 	src_data_115;
output 	src_data_116;
output 	src_data_86;
input 	Selector5;
input 	Selector12;
output 	src_data_80;
input 	Selector6;
input 	Selector13;
output 	src_data_79;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[1]~0_combout ;
wire \arb|grant[0]~1_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~0_combout ;


spw_babasu_altera_merlin_arbitrator_15 arb(
	.nxt_in_ready(nxt_in_ready),
	.nxt_in_ready1(nxt_in_ready1),
	.out_data_4(out_data_4),
	.Equal16(Equal161),
	.Equal161(Equal162),
	.reset(altera_reset_synchronizer_int_chain_out),
	.src16_valid(src16_valid1),
	.src16_valid1(src16_valid3),
	.WideOr1(WideOr11),
	.src_payload_0(src_payload_0),
	.src16_valid2(src16_valid4),
	.grant_1(\arb|grant[1]~0_combout ),
	.packet_in_progress(\packet_in_progress~q ),
	.grant_0(\arb|grant[0]~1_combout ),
	.clk(clk_clk));

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

cyclonev_lcell_comb \src_valid~0 (
	.dataa(!Equal16),
	.datab(!saved_grant_1),
	.datac(!src16_valid2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~0 .extended_lut = "off";
defparam \src_valid~0 .lut_mask = 64'h0101010101010101;
defparam \src_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src_valid~1 (
	.dataa(!out_data_4),
	.datab(!Equal161),
	.datac(!Equal162),
	.datad(!saved_grant_0),
	.datae(!write_addr_data_both_valid),
	.dataf(!src16_valid),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~1 .extended_lut = "off";
defparam \src_valid~1 .lut_mask = 64'h0000000200000000;
defparam \src_valid~1 .shared_arith = "off";

cyclonev_lcell_comb WideOr1(
	.dataa(!out_data_4),
	.datab(!Equal161),
	.datac(!Equal162),
	.datad(!saved_grant_0),
	.datae(!src16_valid3),
	.dataf(!src_valid),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr11),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr1.extended_lut = "off";
defparam WideOr1.lut_mask = 64'hFFFFFFFD00000000;
defparam WideOr1.shared_arith = "off";

cyclonev_lcell_comb \src_data[87] (
	.dataa(!h2f_ARSIZE_1),
	.datab(!h2f_AWSIZE_1),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_87),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[87] .extended_lut = "off";
defparam \src_data[87] .lut_mask = 64'h0537053705370537;
defparam \src_data[87] .shared_arith = "off";

cyclonev_lcell_comb \src_data[88] (
	.dataa(!h2f_ARSIZE_2),
	.datab(!h2f_AWSIZE_2),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_88),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[88] .extended_lut = "off";
defparam \src_data[88] .lut_mask = 64'h0537053705370537;
defparam \src_data[88] .shared_arith = "off";

cyclonev_lcell_comb \src_data[35] (
	.dataa(!h2f_WSTRB_3),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_35),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[35] .extended_lut = "off";
defparam \src_data[35] .lut_mask = 64'h3737373737373737;
defparam \src_data[35] .shared_arith = "off";

cyclonev_lcell_comb \src_data[34] (
	.dataa(!h2f_WSTRB_2),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_34),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[34] .extended_lut = "off";
defparam \src_data[34] .lut_mask = 64'h3737373737373737;
defparam \src_data[34] .shared_arith = "off";

cyclonev_lcell_comb \src_data[33] (
	.dataa(!h2f_WSTRB_1),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_33),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[33] .extended_lut = "off";
defparam \src_data[33] .lut_mask = 64'h3737373737373737;
defparam \src_data[33] .shared_arith = "off";

cyclonev_lcell_comb \src_data[32] (
	.dataa(!h2f_WSTRB_0),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_32),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[32] .extended_lut = "off";
defparam \src_data[32] .lut_mask = 64'h3737373737373737;
defparam \src_data[32] .shared_arith = "off";

cyclonev_lcell_comb \src_payload[0] (
	.dataa(!h2f_WLAST_0),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload[0] .extended_lut = "off";
defparam \src_payload[0] .lut_mask = 64'h3737373737373737;
defparam \src_payload[0] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!h2f_WDATA_0),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h1111111111111111;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[82] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector3),
	.datad(!Selector10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_82),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[82] .extended_lut = "off";
defparam \src_data[82] .lut_mask = 64'h0357035703570357;
defparam \src_data[82] .shared_arith = "off";

cyclonev_lcell_comb \src_data[81] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector4),
	.datad(!Selector11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_81),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[81] .extended_lut = "off";
defparam \src_data[81] .lut_mask = 64'h0357035703570357;
defparam \src_data[81] .shared_arith = "off";

cyclonev_lcell_comb \src_data[105] (
	.dataa(!h2f_ARID_0),
	.datab(!h2f_AWID_0),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_105),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[105] .extended_lut = "off";
defparam \src_data[105] .lut_mask = 64'h0537053705370537;
defparam \src_data[105] .shared_arith = "off";

cyclonev_lcell_comb \src_data[106] (
	.dataa(!h2f_ARID_1),
	.datab(!h2f_AWID_1),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_106),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[106] .extended_lut = "off";
defparam \src_data[106] .lut_mask = 64'h0537053705370537;
defparam \src_data[106] .shared_arith = "off";

cyclonev_lcell_comb \src_data[107] (
	.dataa(!h2f_ARID_2),
	.datab(!h2f_AWID_2),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_107),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[107] .extended_lut = "off";
defparam \src_data[107] .lut_mask = 64'h0537053705370537;
defparam \src_data[107] .shared_arith = "off";

cyclonev_lcell_comb \src_data[108] (
	.dataa(!h2f_ARID_3),
	.datab(!h2f_AWID_3),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_108),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[108] .extended_lut = "off";
defparam \src_data[108] .lut_mask = 64'h0537053705370537;
defparam \src_data[108] .shared_arith = "off";

cyclonev_lcell_comb \src_data[109] (
	.dataa(!h2f_ARID_4),
	.datab(!h2f_AWID_4),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_109),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[109] .extended_lut = "off";
defparam \src_data[109] .lut_mask = 64'h0537053705370537;
defparam \src_data[109] .shared_arith = "off";

cyclonev_lcell_comb \src_data[110] (
	.dataa(!h2f_ARID_5),
	.datab(!h2f_AWID_5),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_110),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[110] .extended_lut = "off";
defparam \src_data[110] .lut_mask = 64'h0537053705370537;
defparam \src_data[110] .shared_arith = "off";

cyclonev_lcell_comb \src_data[111] (
	.dataa(!h2f_ARID_6),
	.datab(!h2f_AWID_6),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_111),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[111] .extended_lut = "off";
defparam \src_data[111] .lut_mask = 64'h0537053705370537;
defparam \src_data[111] .shared_arith = "off";

cyclonev_lcell_comb \src_data[112] (
	.dataa(!h2f_ARID_7),
	.datab(!h2f_AWID_7),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_112),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[112] .extended_lut = "off";
defparam \src_data[112] .lut_mask = 64'h0537053705370537;
defparam \src_data[112] .shared_arith = "off";

cyclonev_lcell_comb \src_data[113] (
	.dataa(!h2f_ARID_8),
	.datab(!h2f_AWID_8),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_113),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[113] .extended_lut = "off";
defparam \src_data[113] .lut_mask = 64'h0537053705370537;
defparam \src_data[113] .shared_arith = "off";

cyclonev_lcell_comb \src_data[114] (
	.dataa(!h2f_ARID_9),
	.datab(!h2f_AWID_9),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_114),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[114] .extended_lut = "off";
defparam \src_data[114] .lut_mask = 64'h0537053705370537;
defparam \src_data[114] .shared_arith = "off";

cyclonev_lcell_comb \src_data[115] (
	.dataa(!h2f_ARID_10),
	.datab(!h2f_AWID_10),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_115),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[115] .extended_lut = "off";
defparam \src_data[115] .lut_mask = 64'h0537053705370537;
defparam \src_data[115] .shared_arith = "off";

cyclonev_lcell_comb \src_data[116] (
	.dataa(!h2f_ARID_11),
	.datab(!h2f_AWID_11),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_116),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[116] .extended_lut = "off";
defparam \src_data[116] .lut_mask = 64'h0537053705370537;
defparam \src_data[116] .shared_arith = "off";

cyclonev_lcell_comb \src_data[86] (
	.dataa(!h2f_ARSIZE_0),
	.datab(!h2f_AWSIZE_0),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_86),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[86] .extended_lut = "off";
defparam \src_data[86] .lut_mask = 64'h0537053705370537;
defparam \src_data[86] .shared_arith = "off";

cyclonev_lcell_comb \src_data[80] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector5),
	.datad(!Selector12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_80),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[80] .extended_lut = "off";
defparam \src_data[80] .lut_mask = 64'h0357035703570357;
defparam \src_data[80] .shared_arith = "off";

cyclonev_lcell_comb \src_data[79] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector6),
	.datad(!Selector13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_79),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[79] .extended_lut = "off";
defparam \src_data[79] .lut_mask = 64'h0357035703570357;
defparam \src_data[79] .shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!\update_grant~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \update_grant~0 (
	.dataa(!nxt_in_ready1),
	.datab(!nxt_in_ready),
	.datac(!src_valid),
	.datad(!src_valid1),
	.datae(!src_payload_0),
	.dataf(!\packet_in_progress~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\update_grant~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \update_grant~0 .extended_lut = "off";
defparam \update_grant~0 .lut_mask = 64'hF000F77700000777;
defparam \update_grant~0 .shared_arith = "off";

endmodule

module spw_babasu_altera_merlin_arbitrator_15 (
	nxt_in_ready,
	nxt_in_ready1,
	out_data_4,
	Equal16,
	Equal161,
	reset,
	src16_valid,
	src16_valid1,
	WideOr1,
	src_payload_0,
	src16_valid2,
	grant_1,
	packet_in_progress,
	grant_0,
	clk)/* synthesis synthesis_greybox=0 */;
input 	nxt_in_ready;
input 	nxt_in_ready1;
input 	out_data_4;
input 	Equal16;
input 	Equal161;
input 	reset;
input 	src16_valid;
input 	src16_valid1;
input 	WideOr1;
input 	src_payload_0;
input 	src16_valid2;
output 	grant_1;
input 	packet_in_progress;
output 	grant_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg[0]~2_combout ;
wire \top_priority_reg[0]~q ;


cyclonev_lcell_comb \grant[1]~0 (
	.dataa(!\top_priority_reg[1]~q ),
	.datab(!\top_priority_reg[0]~q ),
	.datac(!src16_valid),
	.datad(!src16_valid2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[1]~0 .extended_lut = "off";
defparam \grant[1]~0 .lut_mask = 64'h00D500D500D500D5;
defparam \grant[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \grant[0]~1 (
	.dataa(!\top_priority_reg[1]~q ),
	.datab(!\top_priority_reg[0]~q ),
	.datac(!src16_valid),
	.datad(!src16_valid2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[0]~1 .extended_lut = "off";
defparam \grant[0]~1 .lut_mask = 64'h0D0C0D0C0D0C0D0C;
defparam \grant[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~0 (
	.dataa(!out_data_4),
	.datab(!Equal16),
	.datac(!Equal161),
	.datad(!src16_valid1),
	.datae(!src16_valid2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~0 .extended_lut = "off";
defparam \top_priority_reg[0]~0 .lut_mask = 64'hFFFD0000FFFD0000;
defparam \top_priority_reg[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~1 (
	.dataa(!nxt_in_ready1),
	.datab(!nxt_in_ready),
	.datac(!WideOr1),
	.datad(!src_payload_0),
	.datae(!packet_in_progress),
	.dataf(!\top_priority_reg[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~1 .extended_lut = "off";
defparam \top_priority_reg[0]~1 .lut_mask = 64'h0F7F007000000000;
defparam \top_priority_reg[0]~1 .shared_arith = "off";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~1_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

cyclonev_lcell_comb \top_priority_reg[0]~2 (
	.dataa(!grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~2 .extended_lut = "off";
defparam \top_priority_reg[0]~2 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \top_priority_reg[0]~2 .shared_arith = "off";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~1_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

endmodule

module spw_babasu_altera_merlin_arbitrator_16 (
	nxt_in_ready,
	nxt_in_ready1,
	reset,
	src0_valid,
	src0_valid1,
	grant_1,
	src_payload_0,
	packet_in_progress,
	grant_0,
	WideOr1,
	clk)/* synthesis synthesis_greybox=0 */;
input 	nxt_in_ready;
input 	nxt_in_ready1;
input 	reset;
input 	src0_valid;
input 	src0_valid1;
output 	grant_1;
input 	src_payload_0;
input 	packet_in_progress;
output 	grant_0;
input 	WideOr1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg[0]~4_combout ;
wire \top_priority_reg[0]~q ;


cyclonev_lcell_comb \grant[1]~0 (
	.dataa(!\top_priority_reg[1]~q ),
	.datab(!\top_priority_reg[0]~q ),
	.datac(!src0_valid),
	.datad(!src0_valid1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[1]~0 .extended_lut = "off";
defparam \grant[1]~0 .lut_mask = 64'h00D500D500D500D5;
defparam \grant[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \grant[0]~1 (
	.dataa(!\top_priority_reg[1]~q ),
	.datab(!\top_priority_reg[0]~q ),
	.datac(!src0_valid),
	.datad(!src0_valid1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[0]~1 .extended_lut = "off";
defparam \grant[0]~1 .lut_mask = 64'h0D0C0D0C0D0C0D0C;
defparam \grant[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~0 (
	.dataa(!src0_valid1),
	.datab(!src0_valid),
	.datac(!nxt_in_ready),
	.datad(!src_payload_0),
	.datae(!WideOr1),
	.dataf(!nxt_in_ready1),
	.datag(!packet_in_progress),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~0 .extended_lut = "on";
defparam \top_priority_reg[0]~0 .lut_mask = 64'h7070000770700077;
defparam \top_priority_reg[0]~0 .shared_arith = "off";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

cyclonev_lcell_comb \top_priority_reg[0]~4 (
	.dataa(!grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~4 .extended_lut = "off";
defparam \top_priority_reg[0]~4 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \top_priority_reg[0]~4 .shared_arith = "off";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

endmodule

module spw_babasu_spw_babasu_mm_interconnect_0_router (
	h2f_AWADDR_4,
	h2f_AWADDR_5,
	h2f_AWADDR_6,
	h2f_AWADDR_7,
	h2f_AWADDR_8,
	address_burst_8,
	address_burst_7,
	address_burst_6,
	sop_enable,
	out_data_8,
	address_burst_5,
	out_data_5,
	address_burst_4,
	out_data_4,
	out_data_7,
	out_data_6,
	src_data_102,
	Equal5,
	Equal14,
	src_data_100,
	src_data_101,
	Equal16,
	Equal13,
	src_data_103,
	Equal15,
	Equal161,
	Equal9,
	Equal51,
	Equal151,
	Equal141,
	Equal6,
	src_channel,
	Equal152,
	Equal162,
	Equal131,
	Equal142,
	Equal52,
	Equal91,
	src_channel_0,
	Equal2)/* synthesis synthesis_greybox=0 */;
input 	h2f_AWADDR_4;
input 	h2f_AWADDR_5;
input 	h2f_AWADDR_6;
input 	h2f_AWADDR_7;
input 	h2f_AWADDR_8;
input 	address_burst_8;
input 	address_burst_7;
input 	address_burst_6;
input 	sop_enable;
input 	out_data_8;
input 	address_burst_5;
input 	out_data_5;
input 	address_burst_4;
input 	out_data_4;
input 	out_data_7;
input 	out_data_6;
output 	src_data_102;
output 	Equal5;
output 	Equal14;
output 	src_data_100;
output 	src_data_101;
output 	Equal16;
output 	Equal13;
output 	src_data_103;
output 	Equal15;
output 	Equal161;
output 	Equal9;
output 	Equal51;
output 	Equal151;
output 	Equal141;
output 	Equal6;
output 	src_channel;
output 	Equal152;
output 	Equal162;
output 	Equal131;
output 	Equal142;
output 	Equal52;
output 	Equal91;
output 	src_channel_0;
output 	Equal2;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \src_data[102]~0 (
	.dataa(!out_data_8),
	.datab(!out_data_5),
	.datac(!out_data_4),
	.datad(!out_data_7),
	.datae(!out_data_6),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_102),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[102]~0 .extended_lut = "off";
defparam \src_data[102]~0 .lut_mask = 64'h9FFFD7F79FFFD7F7;
defparam \src_data[102]~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal5~0 (
	.dataa(!h2f_AWADDR_6),
	.datab(!h2f_AWADDR_7),
	.datac(!sop_enable),
	.datad(!address_burst_7),
	.datae(!address_burst_6),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal5),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal5~0 .extended_lut = "off";
defparam \Equal5~0 .lut_mask = 64'h40404F4040404F40;
defparam \Equal5~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal14~0 (
	.dataa(!h2f_AWADDR_5),
	.datab(!h2f_AWADDR_8),
	.datac(!sop_enable),
	.datad(!address_burst_8),
	.datae(!address_burst_5),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal14),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal14~0 .extended_lut = "off";
defparam \Equal14~0 .lut_mask = 64'h40404F4040404F40;
defparam \Equal14~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[100]~1 (
	.dataa(!out_data_8),
	.datab(!out_data_5),
	.datac(!out_data_4),
	.datad(!out_data_7),
	.datae(!out_data_6),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_100),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[100]~1 .extended_lut = "off";
defparam \src_data[100]~1 .lut_mask = 64'h4808000048080000;
defparam \src_data[100]~1 .shared_arith = "off";

cyclonev_lcell_comb \src_data[101]~2 (
	.dataa(!out_data_8),
	.datab(!out_data_5),
	.datac(!out_data_4),
	.datad(!out_data_7),
	.datae(!out_data_6),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_101),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[101]~2 .extended_lut = "off";
defparam \src_data[101]~2 .lut_mask = 64'h97FFDFDF97FFDFDF;
defparam \src_data[101]~2 .shared_arith = "off";

cyclonev_lcell_comb \Equal16~0 (
	.dataa(!h2f_AWADDR_6),
	.datab(!h2f_AWADDR_7),
	.datac(!sop_enable),
	.datad(!address_burst_7),
	.datae(!address_burst_6),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal16),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal16~0 .extended_lut = "off";
defparam \Equal16~0 .lut_mask = 64'h8F8080808F808080;
defparam \Equal16~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal13~0 (
	.dataa(!h2f_AWADDR_6),
	.datab(!h2f_AWADDR_7),
	.datac(!sop_enable),
	.datad(!address_burst_7),
	.datae(!address_burst_6),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal13),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal13~0 .extended_lut = "off";
defparam \Equal13~0 .lut_mask = 64'h1010101F1010101F;
defparam \Equal13~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[103]~3 (
	.dataa(!out_data_8),
	.datab(!out_data_5),
	.datac(!out_data_4),
	.datad(!Equal16),
	.datae(!Equal13),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_103),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[103]~3 .extended_lut = "off";
defparam \src_data[103]~3 .lut_mask = 64'h00402A6A00402A6A;
defparam \src_data[103]~3 .shared_arith = "off";

cyclonev_lcell_comb \Equal15~0 (
	.dataa(!h2f_AWADDR_4),
	.datab(!h2f_AWADDR_8),
	.datac(!sop_enable),
	.datad(!address_burst_8),
	.datae(!address_burst_4),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal15),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal15~0 .extended_lut = "off";
defparam \Equal15~0 .lut_mask = 64'h40404F4040404F40;
defparam \Equal15~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal16~1 (
	.dataa(!h2f_AWADDR_5),
	.datab(!h2f_AWADDR_8),
	.datac(!sop_enable),
	.datad(!address_burst_8),
	.datae(!address_burst_5),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal161),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal16~1 .extended_lut = "off";
defparam \Equal16~1 .lut_mask = 64'h202F2020202F2020;
defparam \Equal16~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal9~0 (
	.dataa(!h2f_AWADDR_6),
	.datab(!h2f_AWADDR_7),
	.datac(!sop_enable),
	.datad(!address_burst_7),
	.datae(!address_burst_6),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal9),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal9~0 .extended_lut = "off";
defparam \Equal9~0 .lut_mask = 64'h202F2020202F2020;
defparam \Equal9~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal5~1 (
	.dataa(!h2f_AWADDR_8),
	.datab(!sop_enable),
	.datac(!address_burst_8),
	.datad(!out_data_5),
	.datae(!out_data_4),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal51),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal5~1 .extended_lut = "off";
defparam \Equal5~1 .lut_mask = 64'h0000B8000000B800;
defparam \Equal5~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal15~1 (
	.dataa(!h2f_AWADDR_6),
	.datab(!h2f_AWADDR_7),
	.datac(!sop_enable),
	.datad(!out_data_5),
	.datae(!address_burst_7),
	.dataf(!address_burst_6),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal151),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal15~1 .extended_lut = "off";
defparam \Equal15~1 .lut_mask = 64'h001000100010001F;
defparam \Equal15~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal14~1 (
	.dataa(!h2f_AWADDR_8),
	.datab(!sop_enable),
	.datac(!address_burst_8),
	.datad(!out_data_5),
	.datae(!out_data_4),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal141),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal14~1 .extended_lut = "off";
defparam \Equal14~1 .lut_mask = 64'h00B8000000B80000;
defparam \Equal14~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal6~0 (
	.dataa(!out_data_4),
	.datab(!Equal5),
	.datac(!Equal14),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal6),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal6~0 .extended_lut = "off";
defparam \Equal6~0 .lut_mask = 64'h0202020202020202;
defparam \Equal6~0 .shared_arith = "off";

cyclonev_lcell_comb \src_channel~0 (
	.dataa(!out_data_5),
	.datab(!Equal16),
	.datac(!Equal15),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_channel),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_channel~0 .extended_lut = "off";
defparam \src_channel~0 .lut_mask = 64'h0202020202020202;
defparam \src_channel~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal15~2 (
	.dataa(!out_data_5),
	.datab(!Equal15),
	.datac(!Equal13),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal152),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal15~2 .extended_lut = "off";
defparam \Equal15~2 .lut_mask = 64'h0101010101010101;
defparam \Equal15~2 .shared_arith = "off";

cyclonev_lcell_comb \Equal16~2 (
	.dataa(!out_data_4),
	.datab(!Equal16),
	.datac(!Equal161),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal162),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal16~2 .extended_lut = "off";
defparam \Equal16~2 .lut_mask = 64'h0202020202020202;
defparam \Equal16~2 .shared_arith = "off";

cyclonev_lcell_comb \Equal13~1 (
	.dataa(!out_data_5),
	.datab(!Equal15),
	.datac(!Equal13),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal131),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal13~1 .extended_lut = "off";
defparam \Equal13~1 .lut_mask = 64'h0202020202020202;
defparam \Equal13~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal14~2 (
	.dataa(!out_data_4),
	.datab(!Equal14),
	.datac(!Equal13),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal142),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal14~2 .extended_lut = "off";
defparam \Equal14~2 .lut_mask = 64'h0202020202020202;
defparam \Equal14~2 .shared_arith = "off";

cyclonev_lcell_comb \Equal5~2 (
	.dataa(!out_data_5),
	.datab(!Equal15),
	.datac(!Equal5),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal52),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal5~2 .extended_lut = "off";
defparam \Equal5~2 .lut_mask = 64'h0202020202020202;
defparam \Equal5~2 .shared_arith = "off";

cyclonev_lcell_comb \Equal9~1 (
	.dataa(!out_data_5),
	.datab(!Equal15),
	.datac(!Equal9),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal91),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal9~1 .extended_lut = "off";
defparam \Equal9~1 .lut_mask = 64'h0202020202020202;
defparam \Equal9~1 .shared_arith = "off";

cyclonev_lcell_comb \src_channel[0]~1 (
	.dataa(!out_data_8),
	.datab(!out_data_5),
	.datac(!out_data_4),
	.datad(!out_data_7),
	.datae(!out_data_6),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_channel_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_channel[0]~1 .extended_lut = "off";
defparam \src_channel[0]~1 .lut_mask = 64'h97F7D7D597F7D7D5;
defparam \src_channel[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal2~0 (
	.dataa(!out_data_4),
	.datab(!Equal16),
	.datac(!Equal14),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal2),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~0 .extended_lut = "off";
defparam \Equal2~0 .lut_mask = 64'h0202020202020202;
defparam \Equal2~0 .shared_arith = "off";

endmodule

module spw_babasu_spw_babasu_mm_interconnect_0_router_1 (
	h2f_ARADDR_4,
	h2f_ARADDR_5,
	h2f_ARADDR_6,
	h2f_ARADDR_7,
	h2f_ARADDR_8,
	src_data_102,
	Equal6,
	src_data_100,
	src_data_101,
	src_data_103,
	src_channel,
	src_channel_1,
	Equal15,
	Equal16,
	src_channel_13,
	Equal14,
	Equal3,
	Equal10,
	src_channel_0,
	Equal9,
	Equal4,
	Equal7,
	src_channel_2,
	src_channel1)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARADDR_4;
input 	h2f_ARADDR_5;
input 	h2f_ARADDR_6;
input 	h2f_ARADDR_7;
input 	h2f_ARADDR_8;
output 	src_data_102;
output 	Equal6;
output 	src_data_100;
output 	src_data_101;
output 	src_data_103;
output 	src_channel;
output 	src_channel_1;
output 	Equal15;
output 	Equal16;
output 	src_channel_13;
output 	Equal14;
output 	Equal3;
output 	Equal10;
output 	src_channel_0;
output 	Equal9;
output 	Equal4;
output 	Equal7;
output 	src_channel_2;
output 	src_channel1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \src_data[102]~0 (
	.dataa(!h2f_ARADDR_4),
	.datab(!h2f_ARADDR_5),
	.datac(!h2f_ARADDR_6),
	.datad(!h2f_ARADDR_7),
	.datae(!h2f_ARADDR_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_102),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[102]~0 .extended_lut = "off";
defparam \src_data[102]~0 .lut_mask = 64'hC94B7FFFC94B7FFF;
defparam \src_data[102]~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal6~0 (
	.dataa(!h2f_ARADDR_4),
	.datab(!h2f_ARADDR_5),
	.datac(!h2f_ARADDR_6),
	.datad(!h2f_ARADDR_7),
	.datae(!h2f_ARADDR_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal6),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal6~0 .extended_lut = "off";
defparam \Equal6~0 .lut_mask = 64'h0200000002000000;
defparam \Equal6~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[100]~1 (
	.dataa(!h2f_ARADDR_4),
	.datab(!h2f_ARADDR_5),
	.datac(!h2f_ARADDR_6),
	.datad(!h2f_ARADDR_7),
	.datae(!h2f_ARADDR_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_100),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[100]~1 .extended_lut = "off";
defparam \src_data[100]~1 .lut_mask = 64'h51D8800051D88000;
defparam \src_data[100]~1 .shared_arith = "off";

cyclonev_lcell_comb \src_data[101]~2 (
	.dataa(!h2f_ARADDR_4),
	.datab(!h2f_ARADDR_5),
	.datac(!h2f_ARADDR_6),
	.datad(!h2f_ARADDR_7),
	.datae(!h2f_ARADDR_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_101),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[101]~2 .extended_lut = "off";
defparam \src_data[101]~2 .lut_mask = 64'h85D57FFF85D57FFF;
defparam \src_data[101]~2 .shared_arith = "off";

cyclonev_lcell_comb \src_data[103]~3 (
	.dataa(!h2f_ARADDR_4),
	.datab(!h2f_ARADDR_5),
	.datac(!h2f_ARADDR_6),
	.datad(!h2f_ARADDR_7),
	.datae(!h2f_ARADDR_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_103),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[103]~3 .extended_lut = "off";
defparam \src_data[103]~3 .lut_mask = 64'h013F8000013F8000;
defparam \src_data[103]~3 .shared_arith = "off";

cyclonev_lcell_comb \src_channel~0 (
	.dataa(!h2f_ARADDR_4),
	.datab(!h2f_ARADDR_5),
	.datac(!h2f_ARADDR_6),
	.datad(!h2f_ARADDR_7),
	.datae(!h2f_ARADDR_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_channel),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_channel~0 .extended_lut = "off";
defparam \src_channel~0 .lut_mask = 64'h0080000000800000;
defparam \src_channel~0 .shared_arith = "off";

cyclonev_lcell_comb \src_channel[1]~1 (
	.dataa(!h2f_ARADDR_4),
	.datab(!h2f_ARADDR_5),
	.datac(!h2f_ARADDR_6),
	.datad(!h2f_ARADDR_7),
	.datae(!h2f_ARADDR_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_channel_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_channel[1]~1 .extended_lut = "off";
defparam \src_channel[1]~1 .lut_mask = 64'h4000000040000000;
defparam \src_channel[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal15~0 (
	.dataa(!h2f_ARADDR_4),
	.datab(!h2f_ARADDR_5),
	.datac(!h2f_ARADDR_6),
	.datad(!h2f_ARADDR_7),
	.datae(!h2f_ARADDR_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal15),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal15~0 .extended_lut = "off";
defparam \Equal15~0 .lut_mask = 64'h0001000000010000;
defparam \Equal15~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal16~0 (
	.dataa(!h2f_ARADDR_4),
	.datab(!h2f_ARADDR_5),
	.datac(!h2f_ARADDR_6),
	.datad(!h2f_ARADDR_7),
	.datae(!h2f_ARADDR_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal16),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal16~0 .extended_lut = "off";
defparam \Equal16~0 .lut_mask = 64'h0000800000008000;
defparam \Equal16~0 .shared_arith = "off";

cyclonev_lcell_comb \src_channel[13]~2 (
	.dataa(!h2f_ARADDR_4),
	.datab(!h2f_ARADDR_5),
	.datac(!h2f_ARADDR_6),
	.datad(!h2f_ARADDR_7),
	.datae(!h2f_ARADDR_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_channel_13),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_channel[13]~2 .extended_lut = "off";
defparam \src_channel[13]~2 .lut_mask = 64'h0004000000040000;
defparam \src_channel[13]~2 .shared_arith = "off";

cyclonev_lcell_comb \Equal14~0 (
	.dataa(!h2f_ARADDR_4),
	.datab(!h2f_ARADDR_5),
	.datac(!h2f_ARADDR_6),
	.datad(!h2f_ARADDR_7),
	.datae(!h2f_ARADDR_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal14),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal14~0 .extended_lut = "off";
defparam \Equal14~0 .lut_mask = 64'h0002000000020000;
defparam \Equal14~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal3~0 (
	.dataa(!h2f_ARADDR_4),
	.datab(!h2f_ARADDR_5),
	.datac(!h2f_ARADDR_6),
	.datad(!h2f_ARADDR_7),
	.datae(!h2f_ARADDR_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal3),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~0 .extended_lut = "off";
defparam \Equal3~0 .lut_mask = 64'h1000000010000000;
defparam \Equal3~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal10~0 (
	.dataa(!h2f_ARADDR_4),
	.datab(!h2f_ARADDR_5),
	.datac(!h2f_ARADDR_6),
	.datad(!h2f_ARADDR_7),
	.datae(!h2f_ARADDR_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal10),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal10~0 .extended_lut = "off";
defparam \Equal10~0 .lut_mask = 64'h0020000000200000;
defparam \Equal10~0 .shared_arith = "off";

cyclonev_lcell_comb \src_channel[0]~3 (
	.dataa(!h2f_ARADDR_4),
	.datab(!h2f_ARADDR_5),
	.datac(!h2f_ARADDR_6),
	.datad(!h2f_ARADDR_7),
	.datae(!h2f_ARADDR_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_channel_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_channel[0]~3 .extended_lut = "off";
defparam \src_channel[0]~3 .lut_mask = 64'h80007FFF80007FFF;
defparam \src_channel[0]~3 .shared_arith = "off";

cyclonev_lcell_comb \Equal9~0 (
	.dataa(!h2f_ARADDR_4),
	.datab(!h2f_ARADDR_5),
	.datac(!h2f_ARADDR_6),
	.datad(!h2f_ARADDR_7),
	.datae(!h2f_ARADDR_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal9),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal9~0 .extended_lut = "off";
defparam \Equal9~0 .lut_mask = 64'h0040000000400000;
defparam \Equal9~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal4~0 (
	.dataa(!h2f_ARADDR_4),
	.datab(!h2f_ARADDR_5),
	.datac(!h2f_ARADDR_6),
	.datad(!h2f_ARADDR_7),
	.datae(!h2f_ARADDR_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal4),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal4~0 .extended_lut = "off";
defparam \Equal4~0 .lut_mask = 64'h0800000008000000;
defparam \Equal4~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal7~0 (
	.dataa(!h2f_ARADDR_4),
	.datab(!h2f_ARADDR_5),
	.datac(!h2f_ARADDR_6),
	.datad(!h2f_ARADDR_7),
	.datae(!h2f_ARADDR_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal7),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal7~0 .extended_lut = "off";
defparam \Equal7~0 .lut_mask = 64'h0100000001000000;
defparam \Equal7~0 .shared_arith = "off";

cyclonev_lcell_comb \src_channel[2]~4 (
	.dataa(!h2f_ARADDR_4),
	.datab(!h2f_ARADDR_5),
	.datac(!h2f_ARADDR_6),
	.datad(!h2f_ARADDR_7),
	.datae(!h2f_ARADDR_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_channel_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_channel[2]~4 .extended_lut = "off";
defparam \src_channel[2]~4 .lut_mask = 64'h2000000020000000;
defparam \src_channel[2]~4 .shared_arith = "off";

cyclonev_lcell_comb \src_channel~5 (
	.dataa(!h2f_ARADDR_4),
	.datab(!h2f_ARADDR_5),
	.datac(!h2f_ARADDR_6),
	.datad(!h2f_ARADDR_7),
	.datae(!h2f_ARADDR_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_channel1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_channel~5 .extended_lut = "off";
defparam \src_channel~5 .lut_mask = 64'h0400000004000000;
defparam \src_channel~5 .shared_arith = "off";

endmodule

module spw_babasu_spw_babasu_mm_interconnect_0_rsp_demux (
	h2f_BREADY_0,
	h2f_RREADY_0,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_129_0,
	mem_used_01,
	mem_68_0,
	mem_66_0,
	src0_valid1,
	src1_valid,
	WideOr0)/* synthesis synthesis_greybox=0 */;
input 	h2f_BREADY_0;
input 	h2f_RREADY_0;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	mem_129_0;
input 	mem_used_01;
input 	mem_68_0;
input 	mem_66_0;
output 	src0_valid1;
output 	src1_valid;
output 	WideOr0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb src0_valid(
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_129_0),
	.datad(!mem_used_01),
	.datae(!mem_68_0),
	.dataf(!mem_66_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam src0_valid.extended_lut = "off";
defparam src0_valid.lut_mask = 64'h0000777F00000000;
defparam src0_valid.shared_arith = "off";

cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_129_0),
	.datad(!mem_used_01),
	.datae(!mem_68_0),
	.dataf(!mem_66_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'h8880FFFF88808880;
defparam \src1_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!h2f_BREADY_0),
	.datab(!h2f_RREADY_0),
	.datac(!mem_68_0),
	.datad(!mem_66_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h3533353335333533;
defparam \WideOr0~0 .shared_arith = "off";

endmodule

module spw_babasu_spw_babasu_mm_interconnect_0_rsp_demux_1 (
	h2f_BREADY_0,
	h2f_RREADY_0,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_129_0,
	mem_used_01,
	mem_68_0,
	mem_66_0,
	src0_valid1,
	src1_valid,
	WideOr0)/* synthesis synthesis_greybox=0 */;
input 	h2f_BREADY_0;
input 	h2f_RREADY_0;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	mem_129_0;
input 	mem_used_01;
input 	mem_68_0;
input 	mem_66_0;
output 	src0_valid1;
output 	src1_valid;
output 	WideOr0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb src0_valid(
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_129_0),
	.datad(!mem_used_01),
	.datae(!mem_68_0),
	.dataf(!mem_66_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam src0_valid.extended_lut = "off";
defparam src0_valid.lut_mask = 64'h0000777F00000000;
defparam src0_valid.shared_arith = "off";

cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_129_0),
	.datad(!mem_used_01),
	.datae(!mem_68_0),
	.dataf(!mem_66_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'h8880FFFF88808880;
defparam \src1_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!h2f_BREADY_0),
	.datab(!h2f_RREADY_0),
	.datac(!mem_68_0),
	.datad(!mem_66_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h3533353335333533;
defparam \WideOr0~0 .shared_arith = "off";

endmodule

module spw_babasu_spw_babasu_mm_interconnect_0_rsp_demux_2 (
	h2f_BREADY_0,
	h2f_RREADY_0,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_129_0,
	mem_used_01,
	mem_68_0,
	mem_66_0,
	src0_valid1,
	src1_valid,
	WideOr0)/* synthesis synthesis_greybox=0 */;
input 	h2f_BREADY_0;
input 	h2f_RREADY_0;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	mem_129_0;
input 	mem_used_01;
input 	mem_68_0;
input 	mem_66_0;
output 	src0_valid1;
output 	src1_valid;
output 	WideOr0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb src0_valid(
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_129_0),
	.datad(!mem_used_01),
	.datae(!mem_68_0),
	.dataf(!mem_66_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam src0_valid.extended_lut = "off";
defparam src0_valid.lut_mask = 64'h0000777F00000000;
defparam src0_valid.shared_arith = "off";

cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_129_0),
	.datad(!mem_used_01),
	.datae(!mem_68_0),
	.dataf(!mem_66_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'h8880FFFF88808880;
defparam \src1_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!h2f_BREADY_0),
	.datab(!h2f_RREADY_0),
	.datac(!mem_68_0),
	.datad(!mem_66_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h3533353335333533;
defparam \WideOr0~0 .shared_arith = "off";

endmodule

module spw_babasu_spw_babasu_mm_interconnect_0_rsp_demux_5 (
	h2f_BREADY_0,
	h2f_RREADY_0,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_129_0,
	mem_used_01,
	mem_68_0,
	mem_66_0,
	src0_valid1,
	src1_valid,
	WideOr0)/* synthesis synthesis_greybox=0 */;
input 	h2f_BREADY_0;
input 	h2f_RREADY_0;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	mem_129_0;
input 	mem_used_01;
input 	mem_68_0;
input 	mem_66_0;
output 	src0_valid1;
output 	src1_valid;
output 	WideOr0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb src0_valid(
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_129_0),
	.datad(!mem_used_01),
	.datae(!mem_68_0),
	.dataf(!mem_66_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam src0_valid.extended_lut = "off";
defparam src0_valid.lut_mask = 64'h0000777F00000000;
defparam src0_valid.shared_arith = "off";

cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_129_0),
	.datad(!mem_used_01),
	.datae(!mem_68_0),
	.dataf(!mem_66_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'h8880FFFF88808880;
defparam \src1_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!h2f_BREADY_0),
	.datab(!h2f_RREADY_0),
	.datac(!mem_68_0),
	.datad(!mem_66_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h3533353335333533;
defparam \WideOr0~0 .shared_arith = "off";

endmodule

module spw_babasu_spw_babasu_mm_interconnect_0_rsp_demux_6 (
	h2f_BREADY_0,
	h2f_RREADY_0,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_129_0,
	mem_used_01,
	mem_68_0,
	mem_66_0,
	src0_valid1,
	src1_valid,
	WideOr0)/* synthesis synthesis_greybox=0 */;
input 	h2f_BREADY_0;
input 	h2f_RREADY_0;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	mem_129_0;
input 	mem_used_01;
input 	mem_68_0;
input 	mem_66_0;
output 	src0_valid1;
output 	src1_valid;
output 	WideOr0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb src0_valid(
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_129_0),
	.datad(!mem_used_01),
	.datae(!mem_68_0),
	.dataf(!mem_66_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam src0_valid.extended_lut = "off";
defparam src0_valid.lut_mask = 64'h0000777F00000000;
defparam src0_valid.shared_arith = "off";

cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_129_0),
	.datad(!mem_used_01),
	.datae(!mem_68_0),
	.dataf(!mem_66_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'h8880FFFF88808880;
defparam \src1_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!h2f_BREADY_0),
	.datab(!h2f_RREADY_0),
	.datac(!mem_68_0),
	.datad(!mem_66_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h3533353335333533;
defparam \WideOr0~0 .shared_arith = "off";

endmodule

module spw_babasu_spw_babasu_mm_interconnect_0_rsp_demux_9 (
	h2f_BREADY_0,
	h2f_RREADY_0,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_129_0,
	mem_used_01,
	mem_68_0,
	mem_66_0,
	src0_valid1,
	src1_valid,
	WideOr0)/* synthesis synthesis_greybox=0 */;
input 	h2f_BREADY_0;
input 	h2f_RREADY_0;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	mem_129_0;
input 	mem_used_01;
input 	mem_68_0;
input 	mem_66_0;
output 	src0_valid1;
output 	src1_valid;
output 	WideOr0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb src0_valid(
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_129_0),
	.datad(!mem_used_01),
	.datae(!mem_68_0),
	.dataf(!mem_66_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam src0_valid.extended_lut = "off";
defparam src0_valid.lut_mask = 64'h0000777F00000000;
defparam src0_valid.shared_arith = "off";

cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_129_0),
	.datad(!mem_used_01),
	.datae(!mem_68_0),
	.dataf(!mem_66_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'h8880FFFF88808880;
defparam \src1_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!h2f_BREADY_0),
	.datab(!h2f_RREADY_0),
	.datac(!mem_68_0),
	.datad(!mem_66_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h3533353335333533;
defparam \WideOr0~0 .shared_arith = "off";

endmodule

module spw_babasu_spw_babasu_mm_interconnect_0_rsp_demux_13 (
	h2f_BREADY_0,
	h2f_RREADY_0,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_129_0,
	mem_used_01,
	mem_68_0,
	mem_66_0,
	src0_valid1,
	src1_valid,
	WideOr0)/* synthesis synthesis_greybox=0 */;
input 	h2f_BREADY_0;
input 	h2f_RREADY_0;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	mem_129_0;
input 	mem_used_01;
input 	mem_68_0;
input 	mem_66_0;
output 	src0_valid1;
output 	src1_valid;
output 	WideOr0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb src0_valid(
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_129_0),
	.datad(!mem_used_01),
	.datae(!mem_68_0),
	.dataf(!mem_66_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam src0_valid.extended_lut = "off";
defparam src0_valid.lut_mask = 64'h0000777F00000000;
defparam src0_valid.shared_arith = "off";

cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_129_0),
	.datad(!mem_used_01),
	.datae(!mem_68_0),
	.dataf(!mem_66_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'h8880FFFF88808880;
defparam \src1_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!h2f_BREADY_0),
	.datab(!h2f_RREADY_0),
	.datac(!mem_68_0),
	.datad(!mem_66_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h3533353335333533;
defparam \WideOr0~0 .shared_arith = "off";

endmodule

module spw_babasu_spw_babasu_mm_interconnect_0_rsp_demux_14 (
	h2f_BREADY_0,
	h2f_RREADY_0,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_129_0,
	mem_used_01,
	mem_68_0,
	mem_66_0,
	src0_valid1,
	src1_valid,
	WideOr0)/* synthesis synthesis_greybox=0 */;
input 	h2f_BREADY_0;
input 	h2f_RREADY_0;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	mem_129_0;
input 	mem_used_01;
input 	mem_68_0;
input 	mem_66_0;
output 	src0_valid1;
output 	src1_valid;
output 	WideOr0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb src0_valid(
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_129_0),
	.datad(!mem_used_01),
	.datae(!mem_68_0),
	.dataf(!mem_66_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam src0_valid.extended_lut = "off";
defparam src0_valid.lut_mask = 64'h0000777F00000000;
defparam src0_valid.shared_arith = "off";

cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_129_0),
	.datad(!mem_used_01),
	.datae(!mem_68_0),
	.dataf(!mem_66_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'h8880FFFF88808880;
defparam \src1_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!h2f_BREADY_0),
	.datab(!h2f_RREADY_0),
	.datac(!mem_68_0),
	.datad(!mem_66_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h3533353335333533;
defparam \WideOr0~0 .shared_arith = "off";

endmodule

module spw_babasu_spw_babasu_mm_interconnect_0_rsp_demux_15 (
	h2f_BREADY_0,
	h2f_RREADY_0,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_129_0,
	mem_used_01,
	mem_68_0,
	mem_66_0,
	src0_valid1,
	src1_valid,
	WideOr0)/* synthesis synthesis_greybox=0 */;
input 	h2f_BREADY_0;
input 	h2f_RREADY_0;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	mem_129_0;
input 	mem_used_01;
input 	mem_68_0;
input 	mem_66_0;
output 	src0_valid1;
output 	src1_valid;
output 	WideOr0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb src0_valid(
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_129_0),
	.datad(!mem_used_01),
	.datae(!mem_68_0),
	.dataf(!mem_66_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam src0_valid.extended_lut = "off";
defparam src0_valid.lut_mask = 64'h0000777F00000000;
defparam src0_valid.shared_arith = "off";

cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_129_0),
	.datad(!mem_used_01),
	.datae(!mem_68_0),
	.dataf(!mem_66_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'h8880FFFF88808880;
defparam \src1_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!h2f_BREADY_0),
	.datab(!h2f_RREADY_0),
	.datac(!mem_68_0),
	.datad(!mem_66_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h3533353335333533;
defparam \WideOr0~0 .shared_arith = "off";

endmodule

module spw_babasu_spw_babasu_mm_interconnect_0_rsp_demux_16 (
	h2f_BREADY_0,
	h2f_RREADY_0,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_129_0,
	mem_used_01,
	mem_68_0,
	mem_66_0,
	src0_valid1,
	src1_valid,
	WideOr0)/* synthesis synthesis_greybox=0 */;
input 	h2f_BREADY_0;
input 	h2f_RREADY_0;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	mem_129_0;
input 	mem_used_01;
input 	mem_68_0;
input 	mem_66_0;
output 	src0_valid1;
output 	src1_valid;
output 	WideOr0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb src0_valid(
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_129_0),
	.datad(!mem_used_01),
	.datae(!mem_68_0),
	.dataf(!mem_66_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam src0_valid.extended_lut = "off";
defparam src0_valid.lut_mask = 64'h0000777F00000000;
defparam src0_valid.shared_arith = "off";

cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_129_0),
	.datad(!mem_used_01),
	.datae(!mem_68_0),
	.dataf(!mem_66_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'h8880FFFF88808880;
defparam \src1_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!h2f_BREADY_0),
	.datab(!h2f_RREADY_0),
	.datac(!mem_68_0),
	.datad(!mem_66_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h3533353335333533;
defparam \WideOr0~0 .shared_arith = "off";

endmodule

module spw_babasu_spw_babasu_mm_interconnect_0_rsp_mux (
	mem_66_0,
	src0_valid,
	mem_66_01,
	src0_valid1,
	mem_66_02,
	src0_valid2,
	mem_66_03,
	src0_valid3,
	mem_66_04,
	src0_valid4,
	mem_66_05,
	src0_valid5,
	src0_valid6,
	src0_valid7,
	mem_66_06,
	src0_valid8,
	mem_66_07,
	src0_valid9,
	WideOr11,
	comb,
	mem_130_0,
	last_packet_beat,
	last_packet_beat1,
	comb1,
	mem_130_01,
	last_packet_beat2,
	last_packet_beat3,
	comb2,
	mem_130_02,
	last_packet_beat4,
	last_packet_beat5,
	comb3,
	mem_130_03,
	last_packet_beat6,
	last_packet_beat7,
	comb4,
	mem_130_04,
	last_packet_beat8,
	last_packet_beat9,
	comb5,
	mem_130_05,
	last_packet_beat10,
	last_packet_beat11,
	comb6,
	mem_130_06,
	last_packet_beat12,
	last_packet_beat13,
	mem_130_07,
	mem_130_08,
	comb7,
	mem_130_09,
	last_packet_beat14,
	last_packet_beat15,
	mem_105_0,
	mem_105_01,
	mem_105_02,
	mem_105_03,
	mem_105_04,
	mem_105_05,
	mem_105_06,
	mem_105_07,
	mem_105_08,
	mem_105_09,
	src_data_105,
	mem_106_0,
	mem_106_01,
	mem_106_02,
	mem_106_03,
	mem_106_04,
	mem_106_05,
	mem_106_06,
	mem_106_07,
	mem_106_08,
	mem_106_09,
	src_data_106,
	mem_107_0,
	mem_107_01,
	mem_107_02,
	mem_107_03,
	mem_107_04,
	mem_107_05,
	mem_107_06,
	mem_107_07,
	mem_107_08,
	mem_107_09,
	src_data_107,
	mem_108_0,
	mem_108_01,
	mem_108_02,
	mem_108_03,
	mem_108_04,
	mem_108_05,
	mem_108_06,
	mem_108_07,
	mem_108_08,
	mem_108_09,
	src_data_108,
	mem_109_0,
	mem_109_01,
	mem_109_02,
	mem_109_03,
	mem_109_04,
	mem_109_05,
	mem_109_06,
	mem_109_07,
	mem_109_08,
	mem_109_09,
	src_data_109,
	mem_110_0,
	mem_110_01,
	mem_110_02,
	mem_110_03,
	mem_110_04,
	mem_110_05,
	mem_110_06,
	mem_110_07,
	mem_110_08,
	mem_110_09,
	src_data_110,
	mem_111_0,
	mem_111_01,
	mem_111_02,
	mem_111_03,
	mem_111_04,
	mem_111_05,
	mem_111_06,
	mem_111_07,
	mem_111_08,
	mem_111_09,
	src_data_111,
	mem_112_0,
	mem_112_01,
	mem_112_02,
	mem_112_03,
	mem_112_04,
	mem_112_05,
	mem_112_06,
	mem_112_07,
	mem_112_08,
	mem_112_09,
	src_data_112,
	mem_113_0,
	mem_113_01,
	mem_113_02,
	mem_113_03,
	mem_113_04,
	mem_113_05,
	mem_113_06,
	mem_113_07,
	mem_113_08,
	mem_113_09,
	src_data_113,
	mem_114_0,
	mem_114_01,
	mem_114_02,
	mem_114_03,
	mem_114_04,
	mem_114_05,
	mem_114_06,
	mem_114_07,
	mem_114_08,
	mem_114_09,
	src_data_114,
	mem_115_0,
	mem_115_01,
	mem_115_02,
	mem_115_03,
	mem_115_04,
	mem_115_05,
	mem_115_06,
	mem_115_07,
	mem_115_08,
	mem_115_09,
	src_data_115,
	mem_116_0,
	mem_116_01,
	mem_116_02,
	mem_116_03,
	mem_116_04,
	mem_116_05,
	mem_116_06,
	mem_116_07,
	mem_116_08,
	mem_116_09,
	src_data_116,
	last_packet_beat16,
	last_packet_beat17,
	src_payload,
	src_payload1,
	src_payload_0,
	src_payload_01)/* synthesis synthesis_greybox=0 */;
input 	mem_66_0;
input 	src0_valid;
input 	mem_66_01;
input 	src0_valid1;
input 	mem_66_02;
input 	src0_valid2;
input 	mem_66_03;
input 	src0_valid3;
input 	mem_66_04;
input 	src0_valid4;
input 	mem_66_05;
input 	src0_valid5;
input 	src0_valid6;
input 	src0_valid7;
input 	mem_66_06;
input 	src0_valid8;
input 	mem_66_07;
input 	src0_valid9;
output 	WideOr11;
input 	comb;
input 	mem_130_0;
input 	last_packet_beat;
input 	last_packet_beat1;
input 	comb1;
input 	mem_130_01;
input 	last_packet_beat2;
input 	last_packet_beat3;
input 	comb2;
input 	mem_130_02;
input 	last_packet_beat4;
input 	last_packet_beat5;
input 	comb3;
input 	mem_130_03;
input 	last_packet_beat6;
input 	last_packet_beat7;
input 	comb4;
input 	mem_130_04;
input 	last_packet_beat8;
input 	last_packet_beat9;
input 	comb5;
input 	mem_130_05;
input 	last_packet_beat10;
input 	last_packet_beat11;
input 	comb6;
input 	mem_130_06;
input 	last_packet_beat12;
input 	last_packet_beat13;
input 	mem_130_07;
input 	mem_130_08;
input 	comb7;
input 	mem_130_09;
input 	last_packet_beat14;
input 	last_packet_beat15;
input 	mem_105_0;
input 	mem_105_01;
input 	mem_105_02;
input 	mem_105_03;
input 	mem_105_04;
input 	mem_105_05;
input 	mem_105_06;
input 	mem_105_07;
input 	mem_105_08;
input 	mem_105_09;
output 	src_data_105;
input 	mem_106_0;
input 	mem_106_01;
input 	mem_106_02;
input 	mem_106_03;
input 	mem_106_04;
input 	mem_106_05;
input 	mem_106_06;
input 	mem_106_07;
input 	mem_106_08;
input 	mem_106_09;
output 	src_data_106;
input 	mem_107_0;
input 	mem_107_01;
input 	mem_107_02;
input 	mem_107_03;
input 	mem_107_04;
input 	mem_107_05;
input 	mem_107_06;
input 	mem_107_07;
input 	mem_107_08;
input 	mem_107_09;
output 	src_data_107;
input 	mem_108_0;
input 	mem_108_01;
input 	mem_108_02;
input 	mem_108_03;
input 	mem_108_04;
input 	mem_108_05;
input 	mem_108_06;
input 	mem_108_07;
input 	mem_108_08;
input 	mem_108_09;
output 	src_data_108;
input 	mem_109_0;
input 	mem_109_01;
input 	mem_109_02;
input 	mem_109_03;
input 	mem_109_04;
input 	mem_109_05;
input 	mem_109_06;
input 	mem_109_07;
input 	mem_109_08;
input 	mem_109_09;
output 	src_data_109;
input 	mem_110_0;
input 	mem_110_01;
input 	mem_110_02;
input 	mem_110_03;
input 	mem_110_04;
input 	mem_110_05;
input 	mem_110_06;
input 	mem_110_07;
input 	mem_110_08;
input 	mem_110_09;
output 	src_data_110;
input 	mem_111_0;
input 	mem_111_01;
input 	mem_111_02;
input 	mem_111_03;
input 	mem_111_04;
input 	mem_111_05;
input 	mem_111_06;
input 	mem_111_07;
input 	mem_111_08;
input 	mem_111_09;
output 	src_data_111;
input 	mem_112_0;
input 	mem_112_01;
input 	mem_112_02;
input 	mem_112_03;
input 	mem_112_04;
input 	mem_112_05;
input 	mem_112_06;
input 	mem_112_07;
input 	mem_112_08;
input 	mem_112_09;
output 	src_data_112;
input 	mem_113_0;
input 	mem_113_01;
input 	mem_113_02;
input 	mem_113_03;
input 	mem_113_04;
input 	mem_113_05;
input 	mem_113_06;
input 	mem_113_07;
input 	mem_113_08;
input 	mem_113_09;
output 	src_data_113;
input 	mem_114_0;
input 	mem_114_01;
input 	mem_114_02;
input 	mem_114_03;
input 	mem_114_04;
input 	mem_114_05;
input 	mem_114_06;
input 	mem_114_07;
input 	mem_114_08;
input 	mem_114_09;
output 	src_data_114;
input 	mem_115_0;
input 	mem_115_01;
input 	mem_115_02;
input 	mem_115_03;
input 	mem_115_04;
input 	mem_115_05;
input 	mem_115_06;
input 	mem_115_07;
input 	mem_115_08;
input 	mem_115_09;
output 	src_data_115;
input 	mem_116_0;
input 	mem_116_01;
input 	mem_116_02;
input 	mem_116_03;
input 	mem_116_04;
input 	mem_116_05;
input 	mem_116_06;
input 	mem_116_07;
input 	mem_116_08;
input 	mem_116_09;
output 	src_data_116;
input 	last_packet_beat16;
input 	last_packet_beat17;
output 	src_payload;
output 	src_payload1;
output 	src_payload_0;
output 	src_payload_01;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \WideOr1~0_combout ;
wire \WideOr1~1_combout ;
wire \src_data[105]~0_combout ;
wire \src_data[105]~1_combout ;
wire \src_data[105]~2_combout ;
wire \src_data[105]~3_combout ;
wire \src_data[106]~4_combout ;
wire \src_data[106]~5_combout ;
wire \src_data[106]~6_combout ;
wire \src_data[106]~7_combout ;
wire \src_data[107]~8_combout ;
wire \src_data[107]~9_combout ;
wire \src_data[107]~10_combout ;
wire \src_data[107]~11_combout ;
wire \src_data[108]~12_combout ;
wire \src_data[108]~13_combout ;
wire \src_data[108]~14_combout ;
wire \src_data[108]~15_combout ;
wire \src_data[109]~16_combout ;
wire \src_data[109]~17_combout ;
wire \src_data[109]~18_combout ;
wire \src_data[109]~19_combout ;
wire \src_data[110]~20_combout ;
wire \src_data[110]~21_combout ;
wire \src_data[110]~22_combout ;
wire \src_data[110]~23_combout ;
wire \src_data[111]~24_combout ;
wire \src_data[111]~25_combout ;
wire \src_data[111]~26_combout ;
wire \src_data[111]~27_combout ;
wire \src_data[112]~28_combout ;
wire \src_data[112]~29_combout ;
wire \src_data[112]~30_combout ;
wire \src_data[112]~31_combout ;
wire \src_data[113]~32_combout ;
wire \src_data[113]~33_combout ;
wire \src_data[113]~34_combout ;
wire \src_data[113]~35_combout ;
wire \src_data[114]~36_combout ;
wire \src_data[114]~37_combout ;
wire \src_data[114]~38_combout ;
wire \src_data[114]~39_combout ;
wire \src_data[115]~40_combout ;
wire \src_data[115]~41_combout ;
wire \src_data[115]~42_combout ;
wire \src_data[115]~43_combout ;
wire \src_data[116]~44_combout ;
wire \src_data[116]~45_combout ;
wire \src_data[116]~46_combout ;
wire \src_data[116]~47_combout ;
wire \src_payload~2_combout ;
wire \src_payload~3_combout ;
wire \src_payload~4_combout ;
wire \src_payload~5_combout ;
wire \src_payload~6_combout ;
wire \src_payload~7_combout ;


cyclonev_lcell_comb WideOr1(
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!\WideOr1~0_combout ),
	.datad(!\WideOr1~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr11),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr1.extended_lut = "off";
defparam WideOr1.lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam WideOr1.shared_arith = "off";

cyclonev_lcell_comb \src_data[105] (
	.dataa(!src0_valid8),
	.datab(!src0_valid9),
	.datac(!mem_105_0),
	.datad(!mem_105_01),
	.datae(!\src_data[105]~0_combout ),
	.dataf(!\src_data[105]~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_105),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[105] .extended_lut = "off";
defparam \src_data[105] .lut_mask = 64'hFFFFFFFF0537FFFF;
defparam \src_data[105] .shared_arith = "off";

cyclonev_lcell_comb \src_data[106] (
	.dataa(!src0_valid8),
	.datab(!src0_valid9),
	.datac(!mem_106_0),
	.datad(!mem_106_01),
	.datae(!\src_data[106]~4_combout ),
	.dataf(!\src_data[106]~7_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_106),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[106] .extended_lut = "off";
defparam \src_data[106] .lut_mask = 64'hFFFFFFFF0537FFFF;
defparam \src_data[106] .shared_arith = "off";

cyclonev_lcell_comb \src_data[107] (
	.dataa(!src0_valid8),
	.datab(!src0_valid9),
	.datac(!mem_107_0),
	.datad(!mem_107_01),
	.datae(!\src_data[107]~8_combout ),
	.dataf(!\src_data[107]~11_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_107),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[107] .extended_lut = "off";
defparam \src_data[107] .lut_mask = 64'hFFFFFFFF0537FFFF;
defparam \src_data[107] .shared_arith = "off";

cyclonev_lcell_comb \src_data[108] (
	.dataa(!src0_valid8),
	.datab(!src0_valid9),
	.datac(!mem_108_0),
	.datad(!mem_108_01),
	.datae(!\src_data[108]~12_combout ),
	.dataf(!\src_data[108]~15_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_108),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[108] .extended_lut = "off";
defparam \src_data[108] .lut_mask = 64'hFFFFFFFF0537FFFF;
defparam \src_data[108] .shared_arith = "off";

cyclonev_lcell_comb \src_data[109] (
	.dataa(!src0_valid8),
	.datab(!src0_valid9),
	.datac(!mem_109_0),
	.datad(!mem_109_01),
	.datae(!\src_data[109]~16_combout ),
	.dataf(!\src_data[109]~19_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_109),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[109] .extended_lut = "off";
defparam \src_data[109] .lut_mask = 64'hFFFFFFFF0537FFFF;
defparam \src_data[109] .shared_arith = "off";

cyclonev_lcell_comb \src_data[110] (
	.dataa(!src0_valid8),
	.datab(!src0_valid9),
	.datac(!mem_110_0),
	.datad(!mem_110_01),
	.datae(!\src_data[110]~20_combout ),
	.dataf(!\src_data[110]~23_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_110),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[110] .extended_lut = "off";
defparam \src_data[110] .lut_mask = 64'hFFFFFFFF0537FFFF;
defparam \src_data[110] .shared_arith = "off";

cyclonev_lcell_comb \src_data[111] (
	.dataa(!src0_valid8),
	.datab(!src0_valid9),
	.datac(!mem_111_0),
	.datad(!mem_111_01),
	.datae(!\src_data[111]~24_combout ),
	.dataf(!\src_data[111]~27_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_111),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[111] .extended_lut = "off";
defparam \src_data[111] .lut_mask = 64'hFFFFFFFF0537FFFF;
defparam \src_data[111] .shared_arith = "off";

cyclonev_lcell_comb \src_data[112] (
	.dataa(!src0_valid8),
	.datab(!src0_valid9),
	.datac(!mem_112_0),
	.datad(!mem_112_01),
	.datae(!\src_data[112]~28_combout ),
	.dataf(!\src_data[112]~31_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_112),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[112] .extended_lut = "off";
defparam \src_data[112] .lut_mask = 64'hFFFFFFFF0537FFFF;
defparam \src_data[112] .shared_arith = "off";

cyclonev_lcell_comb \src_data[113] (
	.dataa(!src0_valid8),
	.datab(!src0_valid9),
	.datac(!mem_113_0),
	.datad(!mem_113_01),
	.datae(!\src_data[113]~32_combout ),
	.dataf(!\src_data[113]~35_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_113),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[113] .extended_lut = "off";
defparam \src_data[113] .lut_mask = 64'hFFFFFFFF0537FFFF;
defparam \src_data[113] .shared_arith = "off";

cyclonev_lcell_comb \src_data[114] (
	.dataa(!src0_valid8),
	.datab(!src0_valid9),
	.datac(!mem_114_0),
	.datad(!mem_114_01),
	.datae(!\src_data[114]~36_combout ),
	.dataf(!\src_data[114]~39_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_114),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[114] .extended_lut = "off";
defparam \src_data[114] .lut_mask = 64'hFFFFFFFF0537FFFF;
defparam \src_data[114] .shared_arith = "off";

cyclonev_lcell_comb \src_data[115] (
	.dataa(!src0_valid8),
	.datab(!src0_valid9),
	.datac(!mem_115_0),
	.datad(!mem_115_01),
	.datae(!\src_data[115]~40_combout ),
	.dataf(!\src_data[115]~43_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_115),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[115] .extended_lut = "off";
defparam \src_data[115] .lut_mask = 64'hFFFFFFFF0537FFFF;
defparam \src_data[115] .shared_arith = "off";

cyclonev_lcell_comb \src_data[116] (
	.dataa(!src0_valid8),
	.datab(!src0_valid9),
	.datac(!mem_116_0),
	.datad(!mem_116_01),
	.datae(!\src_data[116]~44_combout ),
	.dataf(!\src_data[116]~47_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_116),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[116] .extended_lut = "off";
defparam \src_data[116] .lut_mask = 64'hFFFFFFFF0537FFFF;
defparam \src_data[116] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!comb7),
	.datab(!mem_66_06),
	.datac(!src0_valid8),
	.datad(!mem_130_09),
	.datae(!last_packet_beat14),
	.dataf(!last_packet_beat15),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h000C000D000D000D;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!comb),
	.datab(!mem_66_07),
	.datac(!src0_valid9),
	.datad(!mem_130_0),
	.datae(!last_packet_beat),
	.dataf(!last_packet_beat1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h000C000D000D000D;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_payload[0]~8 (
	.dataa(!\src_payload~2_combout ),
	.datab(!\src_payload~3_combout ),
	.datac(!\src_payload~4_combout ),
	.datad(!\src_payload~5_combout ),
	.datae(!\src_payload~6_combout ),
	.dataf(!\src_payload~7_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload[0]~8 .extended_lut = "off";
defparam \src_payload[0]~8 .lut_mask = 64'h8000000000000000;
defparam \src_payload[0]~8 .shared_arith = "off";

cyclonev_lcell_comb \src_payload[0]~9 (
	.dataa(!src0_valid6),
	.datab(!src0_valid7),
	.datac(!mem_130_07),
	.datad(!last_packet_beat16),
	.datae(!mem_130_08),
	.dataf(!last_packet_beat17),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload_01),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload[0]~9 .extended_lut = "off";
defparam \src_payload[0]~9 .lut_mask = 64'h0500373305000500;
defparam \src_payload[0]~9 .shared_arith = "off";

cyclonev_lcell_comb \WideOr1~0 (
	.dataa(!src0_valid2),
	.datab(!src0_valid3),
	.datac(!src0_valid4),
	.datad(!src0_valid5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr1~0 .extended_lut = "off";
defparam \WideOr1~0 .lut_mask = 64'h8000800080008000;
defparam \WideOr1~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr1~1 (
	.dataa(!src0_valid6),
	.datab(!src0_valid7),
	.datac(!src0_valid8),
	.datad(!src0_valid9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr1~1 .extended_lut = "off";
defparam \WideOr1~1 .lut_mask = 64'h8000800080008000;
defparam \WideOr1~1 .shared_arith = "off";

cyclonev_lcell_comb \src_data[105]~0 (
	.dataa(!src0_valid6),
	.datab(!src0_valid7),
	.datac(!mem_105_02),
	.datad(!mem_105_03),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[105]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[105]~0 .extended_lut = "off";
defparam \src_data[105]~0 .lut_mask = 64'h0537053705370537;
defparam \src_data[105]~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[105]~1 (
	.dataa(!src0_valid2),
	.datab(!src0_valid3),
	.datac(!mem_105_06),
	.datad(!mem_105_07),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[105]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[105]~1 .extended_lut = "off";
defparam \src_data[105]~1 .lut_mask = 64'h0537053705370537;
defparam \src_data[105]~1 .shared_arith = "off";

cyclonev_lcell_comb \src_data[105]~2 (
	.dataa(!src0_valid5),
	.datab(!src0_valid),
	.datac(!mem_105_08),
	.datad(!mem_105_09),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[105]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[105]~2 .extended_lut = "off";
defparam \src_data[105]~2 .lut_mask = 64'h0537053705370537;
defparam \src_data[105]~2 .shared_arith = "off";

cyclonev_lcell_comb \src_data[105]~3 (
	.dataa(!src0_valid4),
	.datab(!src0_valid1),
	.datac(!mem_105_04),
	.datad(!mem_105_05),
	.datae(!\src_data[105]~1_combout ),
	.dataf(!\src_data[105]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[105]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[105]~3 .extended_lut = "off";
defparam \src_data[105]~3 .lut_mask = 64'hFAC8000000000000;
defparam \src_data[105]~3 .shared_arith = "off";

cyclonev_lcell_comb \src_data[106]~4 (
	.dataa(!src0_valid6),
	.datab(!src0_valid7),
	.datac(!mem_106_02),
	.datad(!mem_106_03),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[106]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[106]~4 .extended_lut = "off";
defparam \src_data[106]~4 .lut_mask = 64'h0537053705370537;
defparam \src_data[106]~4 .shared_arith = "off";

cyclonev_lcell_comb \src_data[106]~5 (
	.dataa(!src0_valid2),
	.datab(!src0_valid3),
	.datac(!mem_106_06),
	.datad(!mem_106_07),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[106]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[106]~5 .extended_lut = "off";
defparam \src_data[106]~5 .lut_mask = 64'h0537053705370537;
defparam \src_data[106]~5 .shared_arith = "off";

cyclonev_lcell_comb \src_data[106]~6 (
	.dataa(!src0_valid5),
	.datab(!src0_valid),
	.datac(!mem_106_08),
	.datad(!mem_106_09),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[106]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[106]~6 .extended_lut = "off";
defparam \src_data[106]~6 .lut_mask = 64'h0537053705370537;
defparam \src_data[106]~6 .shared_arith = "off";

cyclonev_lcell_comb \src_data[106]~7 (
	.dataa(!src0_valid4),
	.datab(!src0_valid1),
	.datac(!mem_106_04),
	.datad(!mem_106_05),
	.datae(!\src_data[106]~5_combout ),
	.dataf(!\src_data[106]~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[106]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[106]~7 .extended_lut = "off";
defparam \src_data[106]~7 .lut_mask = 64'hFAC8000000000000;
defparam \src_data[106]~7 .shared_arith = "off";

cyclonev_lcell_comb \src_data[107]~8 (
	.dataa(!src0_valid6),
	.datab(!src0_valid7),
	.datac(!mem_107_02),
	.datad(!mem_107_03),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[107]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[107]~8 .extended_lut = "off";
defparam \src_data[107]~8 .lut_mask = 64'h0537053705370537;
defparam \src_data[107]~8 .shared_arith = "off";

cyclonev_lcell_comb \src_data[107]~9 (
	.dataa(!src0_valid2),
	.datab(!src0_valid3),
	.datac(!mem_107_06),
	.datad(!mem_107_07),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[107]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[107]~9 .extended_lut = "off";
defparam \src_data[107]~9 .lut_mask = 64'h0537053705370537;
defparam \src_data[107]~9 .shared_arith = "off";

cyclonev_lcell_comb \src_data[107]~10 (
	.dataa(!src0_valid5),
	.datab(!src0_valid),
	.datac(!mem_107_08),
	.datad(!mem_107_09),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[107]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[107]~10 .extended_lut = "off";
defparam \src_data[107]~10 .lut_mask = 64'h0537053705370537;
defparam \src_data[107]~10 .shared_arith = "off";

cyclonev_lcell_comb \src_data[107]~11 (
	.dataa(!src0_valid4),
	.datab(!src0_valid1),
	.datac(!mem_107_04),
	.datad(!mem_107_05),
	.datae(!\src_data[107]~9_combout ),
	.dataf(!\src_data[107]~10_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[107]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[107]~11 .extended_lut = "off";
defparam \src_data[107]~11 .lut_mask = 64'hFAC8000000000000;
defparam \src_data[107]~11 .shared_arith = "off";

cyclonev_lcell_comb \src_data[108]~12 (
	.dataa(!src0_valid6),
	.datab(!src0_valid7),
	.datac(!mem_108_02),
	.datad(!mem_108_03),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[108]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[108]~12 .extended_lut = "off";
defparam \src_data[108]~12 .lut_mask = 64'h0537053705370537;
defparam \src_data[108]~12 .shared_arith = "off";

cyclonev_lcell_comb \src_data[108]~13 (
	.dataa(!src0_valid2),
	.datab(!src0_valid3),
	.datac(!mem_108_06),
	.datad(!mem_108_07),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[108]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[108]~13 .extended_lut = "off";
defparam \src_data[108]~13 .lut_mask = 64'h0537053705370537;
defparam \src_data[108]~13 .shared_arith = "off";

cyclonev_lcell_comb \src_data[108]~14 (
	.dataa(!src0_valid5),
	.datab(!src0_valid),
	.datac(!mem_108_08),
	.datad(!mem_108_09),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[108]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[108]~14 .extended_lut = "off";
defparam \src_data[108]~14 .lut_mask = 64'h0537053705370537;
defparam \src_data[108]~14 .shared_arith = "off";

cyclonev_lcell_comb \src_data[108]~15 (
	.dataa(!src0_valid4),
	.datab(!src0_valid1),
	.datac(!mem_108_04),
	.datad(!mem_108_05),
	.datae(!\src_data[108]~13_combout ),
	.dataf(!\src_data[108]~14_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[108]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[108]~15 .extended_lut = "off";
defparam \src_data[108]~15 .lut_mask = 64'hFAC8000000000000;
defparam \src_data[108]~15 .shared_arith = "off";

cyclonev_lcell_comb \src_data[109]~16 (
	.dataa(!src0_valid6),
	.datab(!src0_valid7),
	.datac(!mem_109_02),
	.datad(!mem_109_03),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[109]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[109]~16 .extended_lut = "off";
defparam \src_data[109]~16 .lut_mask = 64'h0537053705370537;
defparam \src_data[109]~16 .shared_arith = "off";

cyclonev_lcell_comb \src_data[109]~17 (
	.dataa(!src0_valid2),
	.datab(!src0_valid3),
	.datac(!mem_109_06),
	.datad(!mem_109_07),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[109]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[109]~17 .extended_lut = "off";
defparam \src_data[109]~17 .lut_mask = 64'h0537053705370537;
defparam \src_data[109]~17 .shared_arith = "off";

cyclonev_lcell_comb \src_data[109]~18 (
	.dataa(!src0_valid5),
	.datab(!src0_valid),
	.datac(!mem_109_08),
	.datad(!mem_109_09),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[109]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[109]~18 .extended_lut = "off";
defparam \src_data[109]~18 .lut_mask = 64'h0537053705370537;
defparam \src_data[109]~18 .shared_arith = "off";

cyclonev_lcell_comb \src_data[109]~19 (
	.dataa(!src0_valid4),
	.datab(!src0_valid1),
	.datac(!mem_109_04),
	.datad(!mem_109_05),
	.datae(!\src_data[109]~17_combout ),
	.dataf(!\src_data[109]~18_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[109]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[109]~19 .extended_lut = "off";
defparam \src_data[109]~19 .lut_mask = 64'hFAC8000000000000;
defparam \src_data[109]~19 .shared_arith = "off";

cyclonev_lcell_comb \src_data[110]~20 (
	.dataa(!src0_valid6),
	.datab(!src0_valid7),
	.datac(!mem_110_02),
	.datad(!mem_110_03),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[110]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[110]~20 .extended_lut = "off";
defparam \src_data[110]~20 .lut_mask = 64'h0537053705370537;
defparam \src_data[110]~20 .shared_arith = "off";

cyclonev_lcell_comb \src_data[110]~21 (
	.dataa(!src0_valid2),
	.datab(!src0_valid3),
	.datac(!mem_110_06),
	.datad(!mem_110_07),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[110]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[110]~21 .extended_lut = "off";
defparam \src_data[110]~21 .lut_mask = 64'h0537053705370537;
defparam \src_data[110]~21 .shared_arith = "off";

cyclonev_lcell_comb \src_data[110]~22 (
	.dataa(!src0_valid5),
	.datab(!src0_valid),
	.datac(!mem_110_08),
	.datad(!mem_110_09),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[110]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[110]~22 .extended_lut = "off";
defparam \src_data[110]~22 .lut_mask = 64'h0537053705370537;
defparam \src_data[110]~22 .shared_arith = "off";

cyclonev_lcell_comb \src_data[110]~23 (
	.dataa(!src0_valid4),
	.datab(!src0_valid1),
	.datac(!mem_110_04),
	.datad(!mem_110_05),
	.datae(!\src_data[110]~21_combout ),
	.dataf(!\src_data[110]~22_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[110]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[110]~23 .extended_lut = "off";
defparam \src_data[110]~23 .lut_mask = 64'hFAC8000000000000;
defparam \src_data[110]~23 .shared_arith = "off";

cyclonev_lcell_comb \src_data[111]~24 (
	.dataa(!src0_valid6),
	.datab(!src0_valid7),
	.datac(!mem_111_02),
	.datad(!mem_111_03),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[111]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[111]~24 .extended_lut = "off";
defparam \src_data[111]~24 .lut_mask = 64'h0537053705370537;
defparam \src_data[111]~24 .shared_arith = "off";

cyclonev_lcell_comb \src_data[111]~25 (
	.dataa(!src0_valid2),
	.datab(!src0_valid3),
	.datac(!mem_111_06),
	.datad(!mem_111_07),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[111]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[111]~25 .extended_lut = "off";
defparam \src_data[111]~25 .lut_mask = 64'h0537053705370537;
defparam \src_data[111]~25 .shared_arith = "off";

cyclonev_lcell_comb \src_data[111]~26 (
	.dataa(!src0_valid5),
	.datab(!src0_valid),
	.datac(!mem_111_08),
	.datad(!mem_111_09),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[111]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[111]~26 .extended_lut = "off";
defparam \src_data[111]~26 .lut_mask = 64'h0537053705370537;
defparam \src_data[111]~26 .shared_arith = "off";

cyclonev_lcell_comb \src_data[111]~27 (
	.dataa(!src0_valid4),
	.datab(!src0_valid1),
	.datac(!mem_111_04),
	.datad(!mem_111_05),
	.datae(!\src_data[111]~25_combout ),
	.dataf(!\src_data[111]~26_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[111]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[111]~27 .extended_lut = "off";
defparam \src_data[111]~27 .lut_mask = 64'hFAC8000000000000;
defparam \src_data[111]~27 .shared_arith = "off";

cyclonev_lcell_comb \src_data[112]~28 (
	.dataa(!src0_valid6),
	.datab(!src0_valid7),
	.datac(!mem_112_02),
	.datad(!mem_112_03),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[112]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[112]~28 .extended_lut = "off";
defparam \src_data[112]~28 .lut_mask = 64'h0537053705370537;
defparam \src_data[112]~28 .shared_arith = "off";

cyclonev_lcell_comb \src_data[112]~29 (
	.dataa(!src0_valid2),
	.datab(!src0_valid3),
	.datac(!mem_112_06),
	.datad(!mem_112_07),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[112]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[112]~29 .extended_lut = "off";
defparam \src_data[112]~29 .lut_mask = 64'h0537053705370537;
defparam \src_data[112]~29 .shared_arith = "off";

cyclonev_lcell_comb \src_data[112]~30 (
	.dataa(!src0_valid5),
	.datab(!src0_valid),
	.datac(!mem_112_08),
	.datad(!mem_112_09),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[112]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[112]~30 .extended_lut = "off";
defparam \src_data[112]~30 .lut_mask = 64'h0537053705370537;
defparam \src_data[112]~30 .shared_arith = "off";

cyclonev_lcell_comb \src_data[112]~31 (
	.dataa(!src0_valid4),
	.datab(!src0_valid1),
	.datac(!mem_112_04),
	.datad(!mem_112_05),
	.datae(!\src_data[112]~29_combout ),
	.dataf(!\src_data[112]~30_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[112]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[112]~31 .extended_lut = "off";
defparam \src_data[112]~31 .lut_mask = 64'hFAC8000000000000;
defparam \src_data[112]~31 .shared_arith = "off";

cyclonev_lcell_comb \src_data[113]~32 (
	.dataa(!src0_valid6),
	.datab(!src0_valid7),
	.datac(!mem_113_02),
	.datad(!mem_113_03),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[113]~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[113]~32 .extended_lut = "off";
defparam \src_data[113]~32 .lut_mask = 64'h0537053705370537;
defparam \src_data[113]~32 .shared_arith = "off";

cyclonev_lcell_comb \src_data[113]~33 (
	.dataa(!src0_valid2),
	.datab(!src0_valid3),
	.datac(!mem_113_06),
	.datad(!mem_113_07),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[113]~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[113]~33 .extended_lut = "off";
defparam \src_data[113]~33 .lut_mask = 64'h0537053705370537;
defparam \src_data[113]~33 .shared_arith = "off";

cyclonev_lcell_comb \src_data[113]~34 (
	.dataa(!src0_valid5),
	.datab(!src0_valid),
	.datac(!mem_113_08),
	.datad(!mem_113_09),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[113]~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[113]~34 .extended_lut = "off";
defparam \src_data[113]~34 .lut_mask = 64'h0537053705370537;
defparam \src_data[113]~34 .shared_arith = "off";

cyclonev_lcell_comb \src_data[113]~35 (
	.dataa(!src0_valid4),
	.datab(!src0_valid1),
	.datac(!mem_113_04),
	.datad(!mem_113_05),
	.datae(!\src_data[113]~33_combout ),
	.dataf(!\src_data[113]~34_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[113]~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[113]~35 .extended_lut = "off";
defparam \src_data[113]~35 .lut_mask = 64'hFAC8000000000000;
defparam \src_data[113]~35 .shared_arith = "off";

cyclonev_lcell_comb \src_data[114]~36 (
	.dataa(!src0_valid6),
	.datab(!src0_valid7),
	.datac(!mem_114_02),
	.datad(!mem_114_03),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[114]~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[114]~36 .extended_lut = "off";
defparam \src_data[114]~36 .lut_mask = 64'h0537053705370537;
defparam \src_data[114]~36 .shared_arith = "off";

cyclonev_lcell_comb \src_data[114]~37 (
	.dataa(!src0_valid2),
	.datab(!src0_valid3),
	.datac(!mem_114_06),
	.datad(!mem_114_07),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[114]~37_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[114]~37 .extended_lut = "off";
defparam \src_data[114]~37 .lut_mask = 64'h0537053705370537;
defparam \src_data[114]~37 .shared_arith = "off";

cyclonev_lcell_comb \src_data[114]~38 (
	.dataa(!src0_valid5),
	.datab(!src0_valid),
	.datac(!mem_114_08),
	.datad(!mem_114_09),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[114]~38_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[114]~38 .extended_lut = "off";
defparam \src_data[114]~38 .lut_mask = 64'h0537053705370537;
defparam \src_data[114]~38 .shared_arith = "off";

cyclonev_lcell_comb \src_data[114]~39 (
	.dataa(!src0_valid4),
	.datab(!src0_valid1),
	.datac(!mem_114_04),
	.datad(!mem_114_05),
	.datae(!\src_data[114]~37_combout ),
	.dataf(!\src_data[114]~38_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[114]~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[114]~39 .extended_lut = "off";
defparam \src_data[114]~39 .lut_mask = 64'hFAC8000000000000;
defparam \src_data[114]~39 .shared_arith = "off";

cyclonev_lcell_comb \src_data[115]~40 (
	.dataa(!src0_valid6),
	.datab(!src0_valid7),
	.datac(!mem_115_02),
	.datad(!mem_115_03),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[115]~40_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[115]~40 .extended_lut = "off";
defparam \src_data[115]~40 .lut_mask = 64'h0537053705370537;
defparam \src_data[115]~40 .shared_arith = "off";

cyclonev_lcell_comb \src_data[115]~41 (
	.dataa(!src0_valid2),
	.datab(!src0_valid3),
	.datac(!mem_115_06),
	.datad(!mem_115_07),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[115]~41_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[115]~41 .extended_lut = "off";
defparam \src_data[115]~41 .lut_mask = 64'h0537053705370537;
defparam \src_data[115]~41 .shared_arith = "off";

cyclonev_lcell_comb \src_data[115]~42 (
	.dataa(!src0_valid5),
	.datab(!src0_valid),
	.datac(!mem_115_08),
	.datad(!mem_115_09),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[115]~42_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[115]~42 .extended_lut = "off";
defparam \src_data[115]~42 .lut_mask = 64'h0537053705370537;
defparam \src_data[115]~42 .shared_arith = "off";

cyclonev_lcell_comb \src_data[115]~43 (
	.dataa(!src0_valid4),
	.datab(!src0_valid1),
	.datac(!mem_115_04),
	.datad(!mem_115_05),
	.datae(!\src_data[115]~41_combout ),
	.dataf(!\src_data[115]~42_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[115]~43_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[115]~43 .extended_lut = "off";
defparam \src_data[115]~43 .lut_mask = 64'hFAC8000000000000;
defparam \src_data[115]~43 .shared_arith = "off";

cyclonev_lcell_comb \src_data[116]~44 (
	.dataa(!src0_valid6),
	.datab(!src0_valid7),
	.datac(!mem_116_02),
	.datad(!mem_116_03),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[116]~44_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[116]~44 .extended_lut = "off";
defparam \src_data[116]~44 .lut_mask = 64'h0537053705370537;
defparam \src_data[116]~44 .shared_arith = "off";

cyclonev_lcell_comb \src_data[116]~45 (
	.dataa(!src0_valid2),
	.datab(!src0_valid3),
	.datac(!mem_116_06),
	.datad(!mem_116_07),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[116]~45_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[116]~45 .extended_lut = "off";
defparam \src_data[116]~45 .lut_mask = 64'h0537053705370537;
defparam \src_data[116]~45 .shared_arith = "off";

cyclonev_lcell_comb \src_data[116]~46 (
	.dataa(!src0_valid5),
	.datab(!src0_valid),
	.datac(!mem_116_08),
	.datad(!mem_116_09),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[116]~46_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[116]~46 .extended_lut = "off";
defparam \src_data[116]~46 .lut_mask = 64'h0537053705370537;
defparam \src_data[116]~46 .shared_arith = "off";

cyclonev_lcell_comb \src_data[116]~47 (
	.dataa(!src0_valid4),
	.datab(!src0_valid1),
	.datac(!mem_116_04),
	.datad(!mem_116_05),
	.datae(!\src_data[116]~45_combout ),
	.dataf(!\src_data[116]~46_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[116]~47_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[116]~47 .extended_lut = "off";
defparam \src_data[116]~47 .lut_mask = 64'hFAC8000000000000;
defparam \src_data[116]~47 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!comb1),
	.datab(!mem_66_02),
	.datac(!src0_valid2),
	.datad(!mem_130_01),
	.datae(!last_packet_beat2),
	.dataf(!last_packet_beat3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h000C000D000D000D;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~3 (
	.dataa(!comb2),
	.datab(!mem_66_03),
	.datac(!src0_valid3),
	.datad(!mem_130_02),
	.datae(!last_packet_beat4),
	.dataf(!last_packet_beat5),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~3 .extended_lut = "off";
defparam \src_payload~3 .lut_mask = 64'h000C000D000D000D;
defparam \src_payload~3 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~4 (
	.dataa(!comb3),
	.datab(!mem_66_04),
	.datac(!src0_valid4),
	.datad(!mem_130_03),
	.datae(!last_packet_beat6),
	.dataf(!last_packet_beat7),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~4 .extended_lut = "off";
defparam \src_payload~4 .lut_mask = 64'h000C000D000D000D;
defparam \src_payload~4 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~5 (
	.dataa(!comb4),
	.datab(!mem_66_05),
	.datac(!src0_valid5),
	.datad(!mem_130_04),
	.datae(!last_packet_beat8),
	.dataf(!last_packet_beat9),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~5 .extended_lut = "off";
defparam \src_payload~5 .lut_mask = 64'h000C000D000D000D;
defparam \src_payload~5 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~6 (
	.dataa(!comb5),
	.datab(!mem_66_0),
	.datac(!src0_valid),
	.datad(!mem_130_05),
	.datae(!last_packet_beat10),
	.dataf(!last_packet_beat11),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~6 .extended_lut = "off";
defparam \src_payload~6 .lut_mask = 64'h000C000D000D000D;
defparam \src_payload~6 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~7 (
	.dataa(!comb6),
	.datab(!mem_66_01),
	.datac(!src0_valid1),
	.datad(!mem_130_06),
	.datae(!last_packet_beat12),
	.dataf(!last_packet_beat13),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~7 .extended_lut = "off";
defparam \src_payload~7 .lut_mask = 64'h000C000D000D000D;
defparam \src_payload~7 .shared_arith = "off";

endmodule

module spw_babasu_spw_babasu_mm_interconnect_0_rsp_mux_1 (
	read_latency_shift_reg_0,
	mem_used_0,
	mem_66_0,
	read_latency_shift_reg_01,
	mem_used_01,
	mem_66_01,
	read_latency_shift_reg_02,
	mem_used_02,
	mem_66_02,
	read_latency_shift_reg_03,
	mem_used_03,
	mem_66_03,
	read_latency_shift_reg_04,
	mem_used_04,
	mem_66_04,
	mem_66_05,
	read_latency_shift_reg_05,
	mem_used_05,
	mem_66_06,
	mem_66_07,
	mem_66_08,
	read_latency_shift_reg_06,
	mem_used_06,
	mem_66_09,
	comb,
	src1_valid,
	mem_130_0,
	last_packet_beat,
	last_packet_beat1,
	src_payload,
	read_latency_shift_reg_07,
	mem_used_07,
	empty,
	last_packet_beat2,
	mem_130_01,
	read_latency_shift_reg_08,
	mem_used_08,
	empty1,
	mem_66_010,
	mem_used_09,
	last_packet_beat3,
	last_packet_beat4,
	mem_130_02,
	read_latency_shift_reg_09,
	mem_used_010,
	empty2,
	mem_66_011,
	mem_used_011,
	last_packet_beat5,
	last_packet_beat6,
	mem_130_03,
	read_latency_shift_reg_010,
	mem_used_012,
	empty3,
	mem_66_012,
	mem_used_013,
	last_packet_beat7,
	last_packet_beat8,
	mem_130_04,
	mem_130_05,
	read_latency_shift_reg_011,
	mem_used_014,
	empty4,
	mem_66_013,
	mem_used_015,
	last_packet_beat9,
	last_packet_beat10,
	src_payload_0,
	comb1,
	src1_valid1,
	mem_130_06,
	last_packet_beat11,
	last_packet_beat12,
	comb2,
	src1_valid2,
	mem_130_07,
	last_packet_beat13,
	last_packet_beat14,
	comb3,
	src1_valid3,
	mem_130_08,
	last_packet_beat15,
	last_packet_beat16,
	comb4,
	src1_valid4,
	mem_130_09,
	last_packet_beat17,
	last_packet_beat18,
	comb5,
	src1_valid5,
	mem_130_010,
	last_packet_beat19,
	last_packet_beat20,
	mem_130_011,
	read_latency_shift_reg_012,
	mem_used_016,
	empty5,
	mem_66_014,
	mem_used_017,
	last_packet_beat21,
	last_packet_beat22,
	src_payload_01,
	read_latency_shift_reg_013,
	mem_used_018,
	empty6,
	last_packet_beat23,
	comb6,
	src1_valid6,
	mem_130_012,
	last_packet_beat24,
	last_packet_beat25,
	comb7,
	src1_valid7,
	mem_130_013,
	last_packet_beat26,
	last_packet_beat27,
	comb8,
	src1_valid8,
	mem_130_014,
	last_packet_beat28,
	last_packet_beat29,
	comb9,
	src1_valid9,
	mem_130_015,
	last_packet_beat30,
	last_packet_beat31,
	mem_130_016,
	src_payload_02,
	src_payload_03,
	WideOr11,
	mem_105_0,
	mem_105_01,
	mem_105_02,
	mem_105_03,
	mem_105_04,
	mem_105_05,
	mem_105_06,
	mem_105_07,
	mem_105_08,
	mem_105_09,
	mem_106_0,
	mem_106_01,
	mem_106_02,
	mem_106_03,
	mem_106_04,
	mem_106_05,
	mem_106_06,
	mem_106_07,
	mem_106_08,
	mem_106_09,
	mem_107_0,
	mem_107_01,
	mem_107_02,
	mem_107_03,
	mem_107_04,
	mem_107_05,
	mem_107_06,
	mem_107_07,
	mem_107_08,
	mem_107_09,
	mem_108_0,
	mem_108_01,
	mem_108_02,
	mem_108_03,
	mem_108_04,
	mem_108_05,
	mem_108_06,
	mem_108_07,
	mem_108_08,
	mem_108_09,
	mem_109_0,
	mem_109_01,
	mem_109_02,
	mem_109_03,
	mem_109_04,
	mem_109_05,
	mem_109_06,
	mem_109_07,
	mem_109_08,
	mem_109_09,
	mem_110_0,
	mem_110_01,
	mem_110_02,
	mem_110_03,
	mem_110_04,
	mem_110_05,
	mem_110_06,
	mem_110_07,
	mem_110_08,
	mem_110_09,
	mem_111_0,
	mem_111_01,
	mem_111_02,
	mem_111_03,
	mem_111_04,
	mem_111_05,
	mem_111_06,
	mem_111_07,
	mem_111_08,
	mem_111_09,
	mem_112_0,
	mem_112_01,
	mem_112_02,
	mem_112_03,
	mem_112_04,
	mem_112_05,
	mem_112_06,
	mem_112_07,
	mem_112_08,
	mem_112_09,
	mem_113_0,
	mem_113_01,
	mem_113_02,
	mem_113_03,
	mem_113_04,
	mem_113_05,
	mem_113_06,
	mem_113_07,
	mem_113_08,
	mem_113_09,
	mem_114_0,
	mem_114_01,
	mem_114_02,
	mem_114_03,
	mem_114_04,
	mem_114_05,
	mem_114_06,
	mem_114_07,
	mem_114_08,
	mem_114_09,
	mem_115_0,
	mem_115_01,
	mem_115_02,
	mem_115_03,
	mem_115_04,
	mem_115_05,
	mem_115_06,
	mem_115_07,
	mem_115_08,
	mem_115_09,
	mem_116_0,
	mem_116_01,
	mem_116_02,
	mem_116_03,
	mem_116_04,
	mem_116_05,
	mem_116_06,
	mem_116_07,
	mem_116_08,
	mem_116_09,
	av_readdata_pre_0,
	mem_0_0,
	av_readdata_pre_01,
	always4,
	mem_0_01,
	av_readdata_pre_02,
	av_readdata_pre_03,
	mem_0_02,
	av_readdata_pre_04,
	av_readdata_pre_05,
	mem_0_03,
	mem_0_04,
	av_readdata_pre_06,
	mem_0_05,
	av_readdata_pre_07,
	mem_0_06,
	av_readdata_pre_08,
	mem_0_07,
	mem_0_08,
	av_readdata_pre_09,
	mem_0_09,
	av_readdata_pre_010,
	mem_0_010,
	av_readdata_pre_011,
	mem_0_011,
	av_readdata_pre_012,
	mem_0_012,
	av_readdata_pre_013,
	mem_0_013,
	av_readdata_pre_014,
	mem_0_014,
	av_readdata_pre_015,
	always41,
	mem_0_015,
	av_readdata_pre_016,
	always42,
	mem_0_016,
	src_data_0,
	av_readdata_pre_1,
	av_readdata_pre_11,
	mem_1_0,
	mem_1_01,
	mem_1_02,
	av_readdata_pre_12,
	av_readdata_pre_13,
	mem_1_03,
	av_readdata_pre_14,
	mem_1_04,
	av_readdata_pre_15,
	mem_1_05,
	av_readdata_pre_16,
	mem_1_06,
	src_payload1,
	av_readdata_pre_2,
	av_readdata_pre_21,
	mem_2_0,
	mem_2_01,
	mem_2_02,
	av_readdata_pre_22,
	av_readdata_pre_23,
	mem_2_03,
	av_readdata_pre_24,
	mem_2_04,
	av_readdata_pre_25,
	mem_2_05,
	av_readdata_pre_26,
	mem_2_06,
	src_payload2,
	av_readdata_pre_3,
	av_readdata_pre_31,
	mem_3_0,
	mem_3_01,
	mem_3_02,
	av_readdata_pre_32,
	av_readdata_pre_33,
	mem_3_03,
	av_readdata_pre_34,
	mem_3_04,
	av_readdata_pre_35,
	mem_3_05,
	src_payload3,
	av_readdata_pre_4,
	av_readdata_pre_41,
	mem_4_0,
	mem_4_01,
	mem_4_02,
	av_readdata_pre_42,
	av_readdata_pre_43,
	mem_4_03,
	av_readdata_pre_44,
	mem_4_04,
	av_readdata_pre_45,
	mem_4_05,
	src_payload4,
	av_readdata_pre_5,
	av_readdata_pre_51,
	mem_5_0,
	mem_5_01,
	mem_5_02,
	av_readdata_pre_52,
	av_readdata_pre_53,
	mem_5_03,
	av_readdata_pre_54,
	mem_5_04,
	av_readdata_pre_55,
	mem_5_05,
	src_payload5,
	av_readdata_pre_6,
	av_readdata_pre_61,
	mem_6_0,
	mem_6_01,
	mem_6_02,
	av_readdata_pre_62,
	av_readdata_pre_63,
	mem_6_03,
	av_readdata_pre_64,
	mem_6_04,
	av_readdata_pre_65,
	mem_6_05,
	src_payload6,
	av_readdata_pre_7,
	av_readdata_pre_71,
	mem_7_0,
	av_readdata_pre_72,
	mem_7_01,
	mem_7_02,
	mem_7_03,
	av_readdata_pre_73,
	av_readdata_pre_74,
	mem_7_04,
	src_payload7,
	av_readdata_pre_8,
	mem_8_0,
	mem_8_01,
	av_readdata_pre_81,
	mem_8_02,
	av_readdata_pre_82,
	src_payload8,
	mem_9_0,
	av_readdata_pre_9,
	src_payload9,
	mem_10_0,
	av_readdata_pre_10,
	src_payload10,
	mem_105_010,
	mem_105_011,
	mem_105_012,
	mem_105_013,
	mem_105_014,
	mem_105_015,
	mem_105_016,
	src_data_105,
	mem_106_010,
	mem_106_011,
	mem_106_012,
	mem_106_013,
	mem_106_014,
	mem_106_015,
	mem_106_016,
	src_data_106,
	mem_107_010,
	mem_107_011,
	mem_107_012,
	mem_107_013,
	mem_107_014,
	mem_107_015,
	mem_107_016,
	src_data_107,
	mem_108_010,
	mem_108_011,
	mem_108_012,
	mem_108_013,
	mem_108_014,
	mem_108_015,
	mem_108_016,
	src_data_108,
	mem_109_010,
	mem_109_011,
	mem_109_012,
	mem_109_013,
	mem_109_014,
	mem_109_015,
	mem_109_016,
	src_data_109,
	mem_110_010,
	mem_110_011,
	mem_110_012,
	mem_110_013,
	mem_110_014,
	mem_110_015,
	mem_110_016,
	src_data_110,
	mem_111_010,
	mem_111_011,
	mem_111_012,
	mem_111_013,
	mem_111_014,
	mem_111_015,
	mem_111_016,
	src_data_111,
	mem_112_010,
	mem_112_011,
	mem_112_012,
	mem_112_013,
	mem_112_014,
	mem_112_015,
	mem_112_016,
	src_data_112,
	mem_113_010,
	mem_113_011,
	mem_113_012,
	mem_113_013,
	mem_113_014,
	mem_113_015,
	mem_113_016,
	src_data_113,
	mem_114_010,
	mem_114_011,
	mem_114_012,
	mem_114_013,
	mem_114_014,
	mem_114_015,
	mem_114_016,
	src_data_114,
	mem_115_010,
	mem_115_011,
	mem_115_012,
	mem_115_013,
	mem_115_014,
	mem_115_015,
	mem_115_016,
	src_data_115,
	mem_116_010,
	mem_116_011,
	mem_116_012,
	mem_116_013,
	mem_116_014,
	mem_116_015,
	mem_116_016,
	src_data_116)/* synthesis synthesis_greybox=0 */;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	mem_66_0;
input 	read_latency_shift_reg_01;
input 	mem_used_01;
input 	mem_66_01;
input 	read_latency_shift_reg_02;
input 	mem_used_02;
input 	mem_66_02;
input 	read_latency_shift_reg_03;
input 	mem_used_03;
input 	mem_66_03;
input 	read_latency_shift_reg_04;
input 	mem_used_04;
input 	mem_66_04;
input 	mem_66_05;
input 	read_latency_shift_reg_05;
input 	mem_used_05;
input 	mem_66_06;
input 	mem_66_07;
input 	mem_66_08;
input 	read_latency_shift_reg_06;
input 	mem_used_06;
input 	mem_66_09;
input 	comb;
input 	src1_valid;
input 	mem_130_0;
input 	last_packet_beat;
input 	last_packet_beat1;
output 	src_payload;
input 	read_latency_shift_reg_07;
input 	mem_used_07;
input 	empty;
input 	last_packet_beat2;
input 	mem_130_01;
input 	read_latency_shift_reg_08;
input 	mem_used_08;
input 	empty1;
input 	mem_66_010;
input 	mem_used_09;
input 	last_packet_beat3;
input 	last_packet_beat4;
input 	mem_130_02;
input 	read_latency_shift_reg_09;
input 	mem_used_010;
input 	empty2;
input 	mem_66_011;
input 	mem_used_011;
input 	last_packet_beat5;
input 	last_packet_beat6;
input 	mem_130_03;
input 	read_latency_shift_reg_010;
input 	mem_used_012;
input 	empty3;
input 	mem_66_012;
input 	mem_used_013;
input 	last_packet_beat7;
input 	last_packet_beat8;
input 	mem_130_04;
input 	mem_130_05;
input 	read_latency_shift_reg_011;
input 	mem_used_014;
input 	empty4;
input 	mem_66_013;
input 	mem_used_015;
input 	last_packet_beat9;
input 	last_packet_beat10;
output 	src_payload_0;
input 	comb1;
input 	src1_valid1;
input 	mem_130_06;
input 	last_packet_beat11;
input 	last_packet_beat12;
input 	comb2;
input 	src1_valid2;
input 	mem_130_07;
input 	last_packet_beat13;
input 	last_packet_beat14;
input 	comb3;
input 	src1_valid3;
input 	mem_130_08;
input 	last_packet_beat15;
input 	last_packet_beat16;
input 	comb4;
input 	src1_valid4;
input 	mem_130_09;
input 	last_packet_beat17;
input 	last_packet_beat18;
input 	comb5;
input 	src1_valid5;
input 	mem_130_010;
input 	last_packet_beat19;
input 	last_packet_beat20;
input 	mem_130_011;
input 	read_latency_shift_reg_012;
input 	mem_used_016;
input 	empty5;
input 	mem_66_014;
input 	mem_used_017;
input 	last_packet_beat21;
input 	last_packet_beat22;
output 	src_payload_01;
input 	read_latency_shift_reg_013;
input 	mem_used_018;
input 	empty6;
input 	last_packet_beat23;
input 	comb6;
input 	src1_valid6;
input 	mem_130_012;
input 	last_packet_beat24;
input 	last_packet_beat25;
input 	comb7;
input 	src1_valid7;
input 	mem_130_013;
input 	last_packet_beat26;
input 	last_packet_beat27;
input 	comb8;
input 	src1_valid8;
input 	mem_130_014;
input 	last_packet_beat28;
input 	last_packet_beat29;
input 	comb9;
input 	src1_valid9;
input 	mem_130_015;
input 	last_packet_beat30;
input 	last_packet_beat31;
input 	mem_130_016;
output 	src_payload_02;
output 	src_payload_03;
output 	WideOr11;
input 	mem_105_0;
input 	mem_105_01;
input 	mem_105_02;
input 	mem_105_03;
input 	mem_105_04;
input 	mem_105_05;
input 	mem_105_06;
input 	mem_105_07;
input 	mem_105_08;
input 	mem_105_09;
input 	mem_106_0;
input 	mem_106_01;
input 	mem_106_02;
input 	mem_106_03;
input 	mem_106_04;
input 	mem_106_05;
input 	mem_106_06;
input 	mem_106_07;
input 	mem_106_08;
input 	mem_106_09;
input 	mem_107_0;
input 	mem_107_01;
input 	mem_107_02;
input 	mem_107_03;
input 	mem_107_04;
input 	mem_107_05;
input 	mem_107_06;
input 	mem_107_07;
input 	mem_107_08;
input 	mem_107_09;
input 	mem_108_0;
input 	mem_108_01;
input 	mem_108_02;
input 	mem_108_03;
input 	mem_108_04;
input 	mem_108_05;
input 	mem_108_06;
input 	mem_108_07;
input 	mem_108_08;
input 	mem_108_09;
input 	mem_109_0;
input 	mem_109_01;
input 	mem_109_02;
input 	mem_109_03;
input 	mem_109_04;
input 	mem_109_05;
input 	mem_109_06;
input 	mem_109_07;
input 	mem_109_08;
input 	mem_109_09;
input 	mem_110_0;
input 	mem_110_01;
input 	mem_110_02;
input 	mem_110_03;
input 	mem_110_04;
input 	mem_110_05;
input 	mem_110_06;
input 	mem_110_07;
input 	mem_110_08;
input 	mem_110_09;
input 	mem_111_0;
input 	mem_111_01;
input 	mem_111_02;
input 	mem_111_03;
input 	mem_111_04;
input 	mem_111_05;
input 	mem_111_06;
input 	mem_111_07;
input 	mem_111_08;
input 	mem_111_09;
input 	mem_112_0;
input 	mem_112_01;
input 	mem_112_02;
input 	mem_112_03;
input 	mem_112_04;
input 	mem_112_05;
input 	mem_112_06;
input 	mem_112_07;
input 	mem_112_08;
input 	mem_112_09;
input 	mem_113_0;
input 	mem_113_01;
input 	mem_113_02;
input 	mem_113_03;
input 	mem_113_04;
input 	mem_113_05;
input 	mem_113_06;
input 	mem_113_07;
input 	mem_113_08;
input 	mem_113_09;
input 	mem_114_0;
input 	mem_114_01;
input 	mem_114_02;
input 	mem_114_03;
input 	mem_114_04;
input 	mem_114_05;
input 	mem_114_06;
input 	mem_114_07;
input 	mem_114_08;
input 	mem_114_09;
input 	mem_115_0;
input 	mem_115_01;
input 	mem_115_02;
input 	mem_115_03;
input 	mem_115_04;
input 	mem_115_05;
input 	mem_115_06;
input 	mem_115_07;
input 	mem_115_08;
input 	mem_115_09;
input 	mem_116_0;
input 	mem_116_01;
input 	mem_116_02;
input 	mem_116_03;
input 	mem_116_04;
input 	mem_116_05;
input 	mem_116_06;
input 	mem_116_07;
input 	mem_116_08;
input 	mem_116_09;
input 	av_readdata_pre_0;
input 	mem_0_0;
input 	av_readdata_pre_01;
input 	always4;
input 	mem_0_01;
input 	av_readdata_pre_02;
input 	av_readdata_pre_03;
input 	mem_0_02;
input 	av_readdata_pre_04;
input 	av_readdata_pre_05;
input 	mem_0_03;
input 	mem_0_04;
input 	av_readdata_pre_06;
input 	mem_0_05;
input 	av_readdata_pre_07;
input 	mem_0_06;
input 	av_readdata_pre_08;
input 	mem_0_07;
input 	mem_0_08;
input 	av_readdata_pre_09;
input 	mem_0_09;
input 	av_readdata_pre_010;
input 	mem_0_010;
input 	av_readdata_pre_011;
input 	mem_0_011;
input 	av_readdata_pre_012;
input 	mem_0_012;
input 	av_readdata_pre_013;
input 	mem_0_013;
input 	av_readdata_pre_014;
input 	mem_0_014;
input 	av_readdata_pre_015;
input 	always41;
input 	mem_0_015;
input 	av_readdata_pre_016;
input 	always42;
input 	mem_0_016;
output 	src_data_0;
input 	av_readdata_pre_1;
input 	av_readdata_pre_11;
input 	mem_1_0;
input 	mem_1_01;
input 	mem_1_02;
input 	av_readdata_pre_12;
input 	av_readdata_pre_13;
input 	mem_1_03;
input 	av_readdata_pre_14;
input 	mem_1_04;
input 	av_readdata_pre_15;
input 	mem_1_05;
input 	av_readdata_pre_16;
input 	mem_1_06;
output 	src_payload1;
input 	av_readdata_pre_2;
input 	av_readdata_pre_21;
input 	mem_2_0;
input 	mem_2_01;
input 	mem_2_02;
input 	av_readdata_pre_22;
input 	av_readdata_pre_23;
input 	mem_2_03;
input 	av_readdata_pre_24;
input 	mem_2_04;
input 	av_readdata_pre_25;
input 	mem_2_05;
input 	av_readdata_pre_26;
input 	mem_2_06;
output 	src_payload2;
input 	av_readdata_pre_3;
input 	av_readdata_pre_31;
input 	mem_3_0;
input 	mem_3_01;
input 	mem_3_02;
input 	av_readdata_pre_32;
input 	av_readdata_pre_33;
input 	mem_3_03;
input 	av_readdata_pre_34;
input 	mem_3_04;
input 	av_readdata_pre_35;
input 	mem_3_05;
output 	src_payload3;
input 	av_readdata_pre_4;
input 	av_readdata_pre_41;
input 	mem_4_0;
input 	mem_4_01;
input 	mem_4_02;
input 	av_readdata_pre_42;
input 	av_readdata_pre_43;
input 	mem_4_03;
input 	av_readdata_pre_44;
input 	mem_4_04;
input 	av_readdata_pre_45;
input 	mem_4_05;
output 	src_payload4;
input 	av_readdata_pre_5;
input 	av_readdata_pre_51;
input 	mem_5_0;
input 	mem_5_01;
input 	mem_5_02;
input 	av_readdata_pre_52;
input 	av_readdata_pre_53;
input 	mem_5_03;
input 	av_readdata_pre_54;
input 	mem_5_04;
input 	av_readdata_pre_55;
input 	mem_5_05;
output 	src_payload5;
input 	av_readdata_pre_6;
input 	av_readdata_pre_61;
input 	mem_6_0;
input 	mem_6_01;
input 	mem_6_02;
input 	av_readdata_pre_62;
input 	av_readdata_pre_63;
input 	mem_6_03;
input 	av_readdata_pre_64;
input 	mem_6_04;
input 	av_readdata_pre_65;
input 	mem_6_05;
output 	src_payload6;
input 	av_readdata_pre_7;
input 	av_readdata_pre_71;
input 	mem_7_0;
input 	av_readdata_pre_72;
input 	mem_7_01;
input 	mem_7_02;
input 	mem_7_03;
input 	av_readdata_pre_73;
input 	av_readdata_pre_74;
input 	mem_7_04;
output 	src_payload7;
input 	av_readdata_pre_8;
input 	mem_8_0;
input 	mem_8_01;
input 	av_readdata_pre_81;
input 	mem_8_02;
input 	av_readdata_pre_82;
output 	src_payload8;
input 	mem_9_0;
input 	av_readdata_pre_9;
output 	src_payload9;
input 	mem_10_0;
input 	av_readdata_pre_10;
output 	src_payload10;
input 	mem_105_010;
input 	mem_105_011;
input 	mem_105_012;
input 	mem_105_013;
input 	mem_105_014;
input 	mem_105_015;
input 	mem_105_016;
output 	src_data_105;
input 	mem_106_010;
input 	mem_106_011;
input 	mem_106_012;
input 	mem_106_013;
input 	mem_106_014;
input 	mem_106_015;
input 	mem_106_016;
output 	src_data_106;
input 	mem_107_010;
input 	mem_107_011;
input 	mem_107_012;
input 	mem_107_013;
input 	mem_107_014;
input 	mem_107_015;
input 	mem_107_016;
output 	src_data_107;
input 	mem_108_010;
input 	mem_108_011;
input 	mem_108_012;
input 	mem_108_013;
input 	mem_108_014;
input 	mem_108_015;
input 	mem_108_016;
output 	src_data_108;
input 	mem_109_010;
input 	mem_109_011;
input 	mem_109_012;
input 	mem_109_013;
input 	mem_109_014;
input 	mem_109_015;
input 	mem_109_016;
output 	src_data_109;
input 	mem_110_010;
input 	mem_110_011;
input 	mem_110_012;
input 	mem_110_013;
input 	mem_110_014;
input 	mem_110_015;
input 	mem_110_016;
output 	src_data_110;
input 	mem_111_010;
input 	mem_111_011;
input 	mem_111_012;
input 	mem_111_013;
input 	mem_111_014;
input 	mem_111_015;
input 	mem_111_016;
output 	src_data_111;
input 	mem_112_010;
input 	mem_112_011;
input 	mem_112_012;
input 	mem_112_013;
input 	mem_112_014;
input 	mem_112_015;
input 	mem_112_016;
output 	src_data_112;
input 	mem_113_010;
input 	mem_113_011;
input 	mem_113_012;
input 	mem_113_013;
input 	mem_113_014;
input 	mem_113_015;
input 	mem_113_016;
output 	src_data_113;
input 	mem_114_010;
input 	mem_114_011;
input 	mem_114_012;
input 	mem_114_013;
input 	mem_114_014;
input 	mem_114_015;
input 	mem_114_016;
output 	src_data_114;
input 	mem_115_010;
input 	mem_115_011;
input 	mem_115_012;
input 	mem_115_013;
input 	mem_115_014;
input 	mem_115_015;
input 	mem_115_016;
output 	src_data_115;
input 	mem_116_010;
input 	mem_116_011;
input 	mem_116_012;
input 	mem_116_013;
input 	mem_116_014;
input 	mem_116_015;
input 	mem_116_016;
output 	src_data_116;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \src_payload~1_combout ;
wire \src_payload~2_combout ;
wire \src_payload~3_combout ;
wire \src_payload~4_combout ;
wire \src_payload~5_combout ;
wire \src_payload~7_combout ;
wire \src_payload~8_combout ;
wire \src_payload~9_combout ;
wire \src_payload~10_combout ;
wire \src_payload~11_combout ;
wire \src_payload~12_combout ;
wire \src_payload~14_combout ;
wire \src_payload~15_combout ;
wire \src_payload~16_combout ;
wire \src_payload~17_combout ;
wire \src_payload~18_combout ;
wire \WideOr1~0_combout ;
wire \WideOr1~1_combout ;
wire \WideOr1~2_combout ;
wire \src_data[0]~0_combout ;
wire \src_data[0]~1_combout ;
wire \src_payload~20_combout ;
wire \src_payload~21_combout ;
wire \src_data[0]~2_combout ;
wire \src_payload~22_combout ;
wire \src_data[0]~3_combout ;
wire \src_data[0]~4_combout ;
wire \src_data[0]~5_combout ;
wire \src_data[0]~6_combout ;
wire \src_data[0]~7_combout ;
wire \src_data[0]~8_combout ;
wire \src_data[0]~9_combout ;
wire \src_data[0]~10_combout ;
wire \src_data[0]~11_combout ;
wire \src_data[0]~12_combout ;
wire \src_data[0]~13_combout ;
wire \src_data[0]~14_combout ;
wire \src_data[0]~15_combout ;
wire \src_data[0]~16_combout ;
wire \src_data[0]~17_combout ;
wire \src_data[0]~18_combout ;
wire \src_data[0]~19_combout ;
wire \src_payload~23_combout ;
wire \src_payload~24_combout ;
wire \src_payload~25_combout ;
wire \src_payload~26_combout ;
wire \src_payload~27_combout ;
wire \src_payload~28_combout ;
wire \src_payload~29_combout ;
wire \src_payload~31_combout ;
wire \src_payload~32_combout ;
wire \src_payload~33_combout ;
wire \src_payload~34_combout ;
wire \src_payload~35_combout ;
wire \src_payload~36_combout ;
wire \src_payload~37_combout ;
wire \src_payload~39_combout ;
wire \src_payload~40_combout ;
wire \src_payload~41_combout ;
wire \src_payload~42_combout ;
wire \src_payload~43_combout ;
wire \src_payload~44_combout ;
wire \src_payload~46_combout ;
wire \src_payload~47_combout ;
wire \src_payload~48_combout ;
wire \src_payload~49_combout ;
wire \src_payload~50_combout ;
wire \src_payload~51_combout ;
wire \src_payload~53_combout ;
wire \src_payload~54_combout ;
wire \src_payload~55_combout ;
wire \src_payload~56_combout ;
wire \src_payload~57_combout ;
wire \src_payload~58_combout ;
wire \src_payload~60_combout ;
wire \src_payload~61_combout ;
wire \src_payload~62_combout ;
wire \src_payload~63_combout ;
wire \src_payload~64_combout ;
wire \src_payload~65_combout ;
wire \src_payload~67_combout ;
wire \src_payload~68_combout ;
wire \src_payload~69_combout ;
wire \src_payload~70_combout ;
wire \src_payload~71_combout ;
wire \src_payload~73_combout ;
wire \src_payload~74_combout ;
wire \src_data[105]~21_combout ;
wire \src_data[105]~22_combout ;
wire \src_data[105]~23_combout ;
wire \src_data[105]~24_combout ;
wire \src_data[105]~25_combout ;
wire \src_data[105]~26_combout ;
wire \src_data[105]~27_combout ;
wire \src_data[106]~28_combout ;
wire \src_data[106]~29_combout ;
wire \src_data[106]~30_combout ;
wire \src_data[106]~31_combout ;
wire \src_data[106]~32_combout ;
wire \src_data[106]~33_combout ;
wire \src_data[106]~34_combout ;
wire \src_data[107]~35_combout ;
wire \src_data[107]~36_combout ;
wire \src_data[107]~37_combout ;
wire \src_data[107]~38_combout ;
wire \src_data[107]~39_combout ;
wire \src_data[107]~40_combout ;
wire \src_data[107]~41_combout ;
wire \src_data[108]~42_combout ;
wire \src_data[108]~43_combout ;
wire \src_data[108]~44_combout ;
wire \src_data[108]~45_combout ;
wire \src_data[108]~46_combout ;
wire \src_data[108]~47_combout ;
wire \src_data[108]~48_combout ;
wire \src_data[109]~49_combout ;
wire \src_data[109]~50_combout ;
wire \src_data[109]~51_combout ;
wire \src_data[109]~52_combout ;
wire \src_data[109]~53_combout ;
wire \src_data[109]~54_combout ;
wire \src_data[109]~55_combout ;
wire \src_data[110]~56_combout ;
wire \src_data[110]~57_combout ;
wire \src_data[110]~58_combout ;
wire \src_data[110]~59_combout ;
wire \src_data[110]~60_combout ;
wire \src_data[110]~61_combout ;
wire \src_data[110]~62_combout ;
wire \src_data[111]~63_combout ;
wire \src_data[111]~64_combout ;
wire \src_data[111]~65_combout ;
wire \src_data[111]~66_combout ;
wire \src_data[111]~67_combout ;
wire \src_data[111]~68_combout ;
wire \src_data[111]~69_combout ;
wire \src_data[112]~70_combout ;
wire \src_data[112]~71_combout ;
wire \src_data[112]~72_combout ;
wire \src_data[112]~73_combout ;
wire \src_data[112]~74_combout ;
wire \src_data[112]~75_combout ;
wire \src_data[112]~76_combout ;
wire \src_data[113]~77_combout ;
wire \src_data[113]~78_combout ;
wire \src_data[113]~79_combout ;
wire \src_data[113]~80_combout ;
wire \src_data[113]~81_combout ;
wire \src_data[113]~82_combout ;
wire \src_data[113]~83_combout ;
wire \src_data[114]~84_combout ;
wire \src_data[114]~85_combout ;
wire \src_data[114]~86_combout ;
wire \src_data[114]~87_combout ;
wire \src_data[114]~88_combout ;
wire \src_data[114]~89_combout ;
wire \src_data[114]~90_combout ;
wire \src_data[115]~91_combout ;
wire \src_data[115]~92_combout ;
wire \src_data[115]~93_combout ;
wire \src_data[115]~94_combout ;
wire \src_data[115]~95_combout ;
wire \src_data[115]~96_combout ;
wire \src_data[115]~97_combout ;
wire \src_data[116]~98_combout ;
wire \src_data[116]~99_combout ;
wire \src_data[116]~100_combout ;
wire \src_data[116]~101_combout ;
wire \src_data[116]~102_combout ;
wire \src_data[116]~103_combout ;
wire \src_data[116]~104_combout ;


cyclonev_lcell_comb \src_payload~0 (
	.dataa(!comb),
	.datab(!mem_66_09),
	.datac(!src1_valid),
	.datad(!mem_130_0),
	.datae(!last_packet_beat),
	.dataf(!last_packet_beat1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h00C000D000D000D0;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload[0]~6 (
	.dataa(!last_packet_beat2),
	.datab(!\src_payload~1_combout ),
	.datac(!\src_payload~2_combout ),
	.datad(!\src_payload~3_combout ),
	.datae(!\src_payload~4_combout ),
	.dataf(!\src_payload~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload[0]~6 .extended_lut = "off";
defparam \src_payload[0]~6 .lut_mask = 64'hC000400000000000;
defparam \src_payload[0]~6 .shared_arith = "off";

cyclonev_lcell_comb \src_payload[0]~13 (
	.dataa(!\src_payload~7_combout ),
	.datab(!\src_payload~8_combout ),
	.datac(!\src_payload~9_combout ),
	.datad(!\src_payload~10_combout ),
	.datae(!\src_payload~11_combout ),
	.dataf(!\src_payload~12_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload_01),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload[0]~13 .extended_lut = "off";
defparam \src_payload[0]~13 .lut_mask = 64'h8000000000000000;
defparam \src_payload[0]~13 .shared_arith = "off";

cyclonev_lcell_comb \src_payload[0]~19 (
	.dataa(!last_packet_beat23),
	.datab(!\src_payload~14_combout ),
	.datac(!\src_payload~15_combout ),
	.datad(!\src_payload~16_combout ),
	.datae(!\src_payload~17_combout ),
	.dataf(!\src_payload~18_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload_02),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload[0]~19 .extended_lut = "off";
defparam \src_payload[0]~19 .lut_mask = 64'hC000000040000000;
defparam \src_payload[0]~19 .shared_arith = "off";

cyclonev_lcell_comb \src_payload[0] (
	.dataa(!src_payload),
	.datab(!src_payload_0),
	.datac(!src_payload_01),
	.datad(!src_payload_02),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload_03),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload[0] .extended_lut = "off";
defparam \src_payload[0] .lut_mask = 64'hFFFDFFFDFFFDFFFD;
defparam \src_payload[0] .shared_arith = "off";

cyclonev_lcell_comb WideOr1(
	.dataa(!empty1),
	.datab(!src1_valid5),
	.datac(!src1_valid9),
	.datad(!src1_valid),
	.datae(!\WideOr1~1_combout ),
	.dataf(!\WideOr1~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr11),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr1.extended_lut = "off";
defparam WideOr1.lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam WideOr1.shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~20 (
	.dataa(!\src_data[0]~0_combout ),
	.datab(!\src_data[0]~1_combout ),
	.datac(!\src_data[0]~8_combout ),
	.datad(!\src_data[0]~11_combout ),
	.datae(!\src_data[0]~15_combout ),
	.dataf(!\src_data[0]~19_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~20 .extended_lut = "off";
defparam \src_data[0]~20 .lut_mask = 64'hFFFFFFFFFFFFF7FF;
defparam \src_data[0]~20 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~30 (
	.dataa(!\src_payload~20_combout ),
	.datab(!av_readdata_pre_1),
	.datac(!\src_payload~23_combout ),
	.datad(!\src_payload~27_combout ),
	.datae(!\src_payload~29_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~30 .extended_lut = "off";
defparam \src_payload~30 .lut_mask = 64'hFFFFFF1FFFFFFF1F;
defparam \src_payload~30 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~38 (
	.dataa(!\src_payload~20_combout ),
	.datab(!av_readdata_pre_2),
	.datac(!\src_payload~31_combout ),
	.datad(!\src_payload~35_combout ),
	.datae(!\src_payload~37_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~38 .extended_lut = "off";
defparam \src_payload~38 .lut_mask = 64'hFFFFFF1FFFFFFF1F;
defparam \src_payload~38 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~45 (
	.dataa(!\src_payload~22_combout ),
	.datab(!av_readdata_pre_3),
	.datac(!\src_payload~39_combout ),
	.datad(!\src_payload~42_combout ),
	.datae(!\src_payload~44_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~45 .extended_lut = "off";
defparam \src_payload~45 .lut_mask = 64'hFFFFFF1FFFFFFF1F;
defparam \src_payload~45 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~52 (
	.dataa(!\src_payload~22_combout ),
	.datab(!av_readdata_pre_4),
	.datac(!\src_payload~46_combout ),
	.datad(!\src_payload~49_combout ),
	.datae(!\src_payload~51_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~52 .extended_lut = "off";
defparam \src_payload~52 .lut_mask = 64'hFFFFFF1FFFFFFF1F;
defparam \src_payload~52 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~59 (
	.dataa(!\src_payload~22_combout ),
	.datab(!av_readdata_pre_5),
	.datac(!\src_payload~53_combout ),
	.datad(!\src_payload~56_combout ),
	.datae(!\src_payload~58_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~59 .extended_lut = "off";
defparam \src_payload~59 .lut_mask = 64'hFFFFFF1FFFFFFF1F;
defparam \src_payload~59 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~66 (
	.dataa(!\src_payload~22_combout ),
	.datab(!av_readdata_pre_6),
	.datac(!\src_payload~60_combout ),
	.datad(!\src_payload~63_combout ),
	.datae(!\src_payload~65_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~66 .extended_lut = "off";
defparam \src_payload~66 .lut_mask = 64'hFFFFFF1FFFFFFF1F;
defparam \src_payload~66 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~72 (
	.dataa(!\src_payload~22_combout ),
	.datab(!av_readdata_pre_7),
	.datac(!\src_payload~67_combout ),
	.datad(!\src_payload~68_combout ),
	.datae(!\src_payload~71_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~72 .extended_lut = "off";
defparam \src_payload~72 .lut_mask = 64'hFFFF1FFFFFFF1FFF;
defparam \src_payload~72 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~75 (
	.dataa(!src1_valid4),
	.datab(!always41),
	.datac(!av_readdata_pre_8),
	.datad(!mem_8_0),
	.datae(!\src_payload~74_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~75 .extended_lut = "off";
defparam \src_payload~75 .lut_mask = 64'hFFFF028AFFFF028A;
defparam \src_payload~75 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~76 (
	.dataa(!read_latency_shift_reg_013),
	.datab(!mem_used_018),
	.datac(!mem_9_0),
	.datad(!av_readdata_pre_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~76 .extended_lut = "off";
defparam \src_payload~76 .lut_mask = 64'h0347034703470347;
defparam \src_payload~76 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~77 (
	.dataa(!read_latency_shift_reg_013),
	.datab(!mem_used_018),
	.datac(!mem_10_0),
	.datad(!av_readdata_pre_10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload10),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~77 .extended_lut = "off";
defparam \src_payload~77 .lut_mask = 64'h0347034703470347;
defparam \src_payload~77 .shared_arith = "off";

cyclonev_lcell_comb \src_data[105] (
	.dataa(!empty1),
	.datab(!mem_105_010),
	.datac(!\src_data[105]~24_combout ),
	.datad(!\src_data[105]~25_combout ),
	.datae(!\src_data[105]~26_combout ),
	.dataf(!\src_data[105]~27_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_105),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[105] .extended_lut = "off";
defparam \src_data[105] .lut_mask = 64'hFFFFFFFFFFFFFFF2;
defparam \src_data[105] .shared_arith = "off";

cyclonev_lcell_comb \src_data[106] (
	.dataa(!empty1),
	.datab(!mem_106_010),
	.datac(!\src_data[106]~31_combout ),
	.datad(!\src_data[106]~32_combout ),
	.datae(!\src_data[106]~33_combout ),
	.dataf(!\src_data[106]~34_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_106),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[106] .extended_lut = "off";
defparam \src_data[106] .lut_mask = 64'hFFFFFFFFFFFFFFF2;
defparam \src_data[106] .shared_arith = "off";

cyclonev_lcell_comb \src_data[107] (
	.dataa(!empty1),
	.datab(!mem_107_010),
	.datac(!\src_data[107]~38_combout ),
	.datad(!\src_data[107]~39_combout ),
	.datae(!\src_data[107]~40_combout ),
	.dataf(!\src_data[107]~41_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_107),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[107] .extended_lut = "off";
defparam \src_data[107] .lut_mask = 64'hFFFFFFFFFFFFFFF2;
defparam \src_data[107] .shared_arith = "off";

cyclonev_lcell_comb \src_data[108] (
	.dataa(!empty1),
	.datab(!mem_108_010),
	.datac(!\src_data[108]~45_combout ),
	.datad(!\src_data[108]~46_combout ),
	.datae(!\src_data[108]~47_combout ),
	.dataf(!\src_data[108]~48_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_108),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[108] .extended_lut = "off";
defparam \src_data[108] .lut_mask = 64'hFFFFFFFFFFFFFFF2;
defparam \src_data[108] .shared_arith = "off";

cyclonev_lcell_comb \src_data[109] (
	.dataa(!empty1),
	.datab(!mem_109_010),
	.datac(!\src_data[109]~52_combout ),
	.datad(!\src_data[109]~53_combout ),
	.datae(!\src_data[109]~54_combout ),
	.dataf(!\src_data[109]~55_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_109),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[109] .extended_lut = "off";
defparam \src_data[109] .lut_mask = 64'hFFFFFFFFFFFFFFF2;
defparam \src_data[109] .shared_arith = "off";

cyclonev_lcell_comb \src_data[110] (
	.dataa(!empty1),
	.datab(!mem_110_010),
	.datac(!\src_data[110]~59_combout ),
	.datad(!\src_data[110]~60_combout ),
	.datae(!\src_data[110]~61_combout ),
	.dataf(!\src_data[110]~62_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_110),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[110] .extended_lut = "off";
defparam \src_data[110] .lut_mask = 64'hFFFFFFFFFFFFFFF2;
defparam \src_data[110] .shared_arith = "off";

cyclonev_lcell_comb \src_data[111] (
	.dataa(!empty1),
	.datab(!mem_111_010),
	.datac(!\src_data[111]~66_combout ),
	.datad(!\src_data[111]~67_combout ),
	.datae(!\src_data[111]~68_combout ),
	.dataf(!\src_data[111]~69_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_111),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[111] .extended_lut = "off";
defparam \src_data[111] .lut_mask = 64'hFFFFFFFFFFFFFFF2;
defparam \src_data[111] .shared_arith = "off";

cyclonev_lcell_comb \src_data[112] (
	.dataa(!empty1),
	.datab(!mem_112_010),
	.datac(!\src_data[112]~73_combout ),
	.datad(!\src_data[112]~74_combout ),
	.datae(!\src_data[112]~75_combout ),
	.dataf(!\src_data[112]~76_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_112),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[112] .extended_lut = "off";
defparam \src_data[112] .lut_mask = 64'hFFFFFFFFFFFFFFF2;
defparam \src_data[112] .shared_arith = "off";

cyclonev_lcell_comb \src_data[113] (
	.dataa(!empty1),
	.datab(!mem_113_010),
	.datac(!\src_data[113]~80_combout ),
	.datad(!\src_data[113]~81_combout ),
	.datae(!\src_data[113]~82_combout ),
	.dataf(!\src_data[113]~83_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_113),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[113] .extended_lut = "off";
defparam \src_data[113] .lut_mask = 64'hFFFFFFFFFFFFFFF2;
defparam \src_data[113] .shared_arith = "off";

cyclonev_lcell_comb \src_data[114] (
	.dataa(!empty1),
	.datab(!mem_114_010),
	.datac(!\src_data[114]~87_combout ),
	.datad(!\src_data[114]~88_combout ),
	.datae(!\src_data[114]~89_combout ),
	.dataf(!\src_data[114]~90_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_114),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[114] .extended_lut = "off";
defparam \src_data[114] .lut_mask = 64'hFFFFFFFFFFFFFFF2;
defparam \src_data[114] .shared_arith = "off";

cyclonev_lcell_comb \src_data[115] (
	.dataa(!empty1),
	.datab(!mem_115_010),
	.datac(!\src_data[115]~94_combout ),
	.datad(!\src_data[115]~95_combout ),
	.datae(!\src_data[115]~96_combout ),
	.dataf(!\src_data[115]~97_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_115),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[115] .extended_lut = "off";
defparam \src_data[115] .lut_mask = 64'hFFFFFFFFFFFFFFF2;
defparam \src_data[115] .shared_arith = "off";

cyclonev_lcell_comb \src_data[116] (
	.dataa(!empty1),
	.datab(!mem_116_010),
	.datac(!\src_data[116]~101_combout ),
	.datad(!\src_data[116]~102_combout ),
	.datae(!\src_data[116]~103_combout ),
	.dataf(!\src_data[116]~104_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_116),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[116] .extended_lut = "off";
defparam \src_data[116] .lut_mask = 64'hFFFFFFFFFFFFFFF2;
defparam \src_data[116] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!mem_130_01),
	.datab(!empty1),
	.datac(!mem_66_010),
	.datad(!mem_used_09),
	.datae(!last_packet_beat3),
	.dataf(!last_packet_beat4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h4040404440444044;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!mem_130_02),
	.datab(!empty2),
	.datac(!mem_66_011),
	.datad(!mem_used_011),
	.datae(!last_packet_beat5),
	.dataf(!last_packet_beat6),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h4040404440444044;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~3 (
	.dataa(!mem_130_03),
	.datab(!empty3),
	.datac(!mem_66_012),
	.datad(!mem_used_013),
	.datae(!last_packet_beat7),
	.dataf(!last_packet_beat8),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~3 .extended_lut = "off";
defparam \src_payload~3 .lut_mask = 64'h4040404440444044;
defparam \src_payload~3 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~4 (
	.dataa(!mem_130_04),
	.datab(!read_latency_shift_reg_07),
	.datac(!mem_used_07),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~4 .extended_lut = "off";
defparam \src_payload~4 .lut_mask = 64'h1515151515151515;
defparam \src_payload~4 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~5 (
	.dataa(!mem_130_05),
	.datab(!empty4),
	.datac(!mem_66_013),
	.datad(!mem_used_015),
	.datae(!last_packet_beat9),
	.dataf(!last_packet_beat10),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~5 .extended_lut = "off";
defparam \src_payload~5 .lut_mask = 64'h4040404440444044;
defparam \src_payload~5 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~7 (
	.dataa(!comb1),
	.datab(!mem_66_02),
	.datac(!src1_valid1),
	.datad(!mem_130_06),
	.datae(!last_packet_beat11),
	.dataf(!last_packet_beat12),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~7 .extended_lut = "off";
defparam \src_payload~7 .lut_mask = 64'h00C000D000D000D0;
defparam \src_payload~7 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~8 (
	.dataa(!comb2),
	.datab(!mem_66_03),
	.datac(!src1_valid2),
	.datad(!mem_130_07),
	.datae(!last_packet_beat13),
	.dataf(!last_packet_beat14),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~8 .extended_lut = "off";
defparam \src_payload~8 .lut_mask = 64'h00C000D000D000D0;
defparam \src_payload~8 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~9 (
	.dataa(!comb3),
	.datab(!mem_66_04),
	.datac(!src1_valid3),
	.datad(!mem_130_08),
	.datae(!last_packet_beat15),
	.dataf(!last_packet_beat16),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~9 .extended_lut = "off";
defparam \src_payload~9 .lut_mask = 64'h00C000D000D000D0;
defparam \src_payload~9 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~10 (
	.dataa(!comb4),
	.datab(!mem_66_05),
	.datac(!src1_valid4),
	.datad(!mem_130_09),
	.datae(!last_packet_beat17),
	.dataf(!last_packet_beat18),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~10 .extended_lut = "off";
defparam \src_payload~10 .lut_mask = 64'h00C000D000D000D0;
defparam \src_payload~10 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~11 (
	.dataa(!comb5),
	.datab(!mem_66_0),
	.datac(!src1_valid5),
	.datad(!mem_130_010),
	.datae(!last_packet_beat19),
	.dataf(!last_packet_beat20),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~11 .extended_lut = "off";
defparam \src_payload~11 .lut_mask = 64'h00C000D000D000D0;
defparam \src_payload~11 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~12 (
	.dataa(!mem_130_011),
	.datab(!empty5),
	.datac(!mem_66_014),
	.datad(!mem_used_017),
	.datae(!last_packet_beat21),
	.dataf(!last_packet_beat22),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~12 .extended_lut = "off";
defparam \src_payload~12 .lut_mask = 64'h4040404440444044;
defparam \src_payload~12 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~14 (
	.dataa(!comb6),
	.datab(!mem_66_01),
	.datac(!src1_valid6),
	.datad(!mem_130_012),
	.datae(!last_packet_beat24),
	.dataf(!last_packet_beat25),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~14 .extended_lut = "off";
defparam \src_payload~14 .lut_mask = 64'h00C000D000D000D0;
defparam \src_payload~14 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~15 (
	.dataa(!comb7),
	.datab(!mem_66_06),
	.datac(!src1_valid7),
	.datad(!mem_130_013),
	.datae(!last_packet_beat26),
	.dataf(!last_packet_beat27),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~15 .extended_lut = "off";
defparam \src_payload~15 .lut_mask = 64'h00C000D000D000D0;
defparam \src_payload~15 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~16 (
	.dataa(!comb8),
	.datab(!mem_66_07),
	.datac(!src1_valid8),
	.datad(!mem_130_014),
	.datae(!last_packet_beat28),
	.dataf(!last_packet_beat29),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~16 .extended_lut = "off";
defparam \src_payload~16 .lut_mask = 64'h00C000D000D000D0;
defparam \src_payload~16 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~17 (
	.dataa(!comb9),
	.datab(!mem_66_08),
	.datac(!src1_valid9),
	.datad(!mem_130_015),
	.datae(!last_packet_beat30),
	.dataf(!last_packet_beat31),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~17 .extended_lut = "off";
defparam \src_payload~17 .lut_mask = 64'h00C000D000D000D0;
defparam \src_payload~17 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~18 (
	.dataa(!mem_130_016),
	.datab(!read_latency_shift_reg_013),
	.datac(!mem_used_018),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~18 .extended_lut = "off";
defparam \src_payload~18 .lut_mask = 64'h1515151515151515;
defparam \src_payload~18 .shared_arith = "off";

cyclonev_lcell_comb \WideOr1~0 (
	.dataa(!read_latency_shift_reg_012),
	.datab(!mem_used_016),
	.datac(!read_latency_shift_reg_013),
	.datad(!mem_used_018),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr1~0 .extended_lut = "off";
defparam \WideOr1~0 .lut_mask = 64'h8000800080008000;
defparam \WideOr1~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr1~1 (
	.dataa(!empty),
	.datab(!src1_valid1),
	.datac(!src1_valid2),
	.datad(!src1_valid3),
	.datae(!src1_valid4),
	.dataf(!\WideOr1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr1~1 .extended_lut = "off";
defparam \WideOr1~1 .lut_mask = 64'h0000000000000001;
defparam \WideOr1~1 .shared_arith = "off";

cyclonev_lcell_comb \WideOr1~2 (
	.dataa(!empty4),
	.datab(!empty3),
	.datac(!empty2),
	.datad(!src1_valid6),
	.datae(!src1_valid7),
	.dataf(!src1_valid8),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr1~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr1~2 .extended_lut = "off";
defparam \WideOr1~2 .lut_mask = 64'h0000000000000001;
defparam \WideOr1~2 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~0 (
	.dataa(!read_latency_shift_reg_04),
	.datab(!mem_used_04),
	.datac(!src1_valid3),
	.datad(!av_readdata_pre_0),
	.datae(!mem_0_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~0 .extended_lut = "off";
defparam \src_data[0]~0 .lut_mask = 64'h0040B0F00040B0F0;
defparam \src_data[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~1 (
	.dataa(!src1_valid9),
	.datab(!av_readdata_pre_01),
	.datac(!always4),
	.datad(!mem_0_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~1 .extended_lut = "off";
defparam \src_data[0]~1 .lut_mask = 64'h02A202A202A202A2;
defparam \src_data[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~20 (
	.dataa(!read_latency_shift_reg_012),
	.datab(!mem_used_016),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~20 .extended_lut = "off";
defparam \src_payload~20 .lut_mask = 64'h4444444444444444;
defparam \src_payload~20 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~21 (
	.dataa(!read_latency_shift_reg_011),
	.datab(!mem_used_014),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~21 .extended_lut = "off";
defparam \src_payload~21 .lut_mask = 64'h4444444444444444;
defparam \src_payload~21 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~2 (
	.dataa(!mem_used_07),
	.datab(!av_readdata_pre_03),
	.datac(!\src_payload~21_combout ),
	.datad(!mem_0_02),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~2 .extended_lut = "off";
defparam \src_data[0]~2 .lut_mask = 64'h0357035703570357;
defparam \src_data[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~22 (
	.dataa(!read_latency_shift_reg_013),
	.datab(!mem_used_018),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~22 .extended_lut = "off";
defparam \src_payload~22 .lut_mask = 64'h4444444444444444;
defparam \src_payload~22 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~3 (
	.dataa(!read_latency_shift_reg_07),
	.datab(!mem_used_07),
	.datac(!av_readdata_pre_04),
	.datad(!av_readdata_pre_05),
	.datae(!\src_payload~22_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~3 .extended_lut = "off";
defparam \src_data[0]~3 .lut_mask = 64'h040404FF040404FF;
defparam \src_data[0]~3 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~4 (
	.dataa(!mem_used_014),
	.datab(!read_latency_shift_reg_08),
	.datac(!mem_used_08),
	.datad(!mem_0_04),
	.datae(!av_readdata_pre_06),
	.dataf(!mem_0_05),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~4 .extended_lut = "off";
defparam \src_data[0]~4 .lut_mask = 64'hFFF0CFC0AAA08A80;
defparam \src_data[0]~4 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~5 (
	.dataa(!read_latency_shift_reg_09),
	.datab(!mem_used_010),
	.datac(!av_readdata_pre_07),
	.datad(!mem_0_06),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[0]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~5 .extended_lut = "off";
defparam \src_data[0]~5 .lut_mask = 64'h0437043704370437;
defparam \src_data[0]~5 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~6 (
	.dataa(!mem_used_016),
	.datab(!read_latency_shift_reg_010),
	.datac(!mem_used_012),
	.datad(!av_readdata_pre_08),
	.datae(!mem_0_07),
	.dataf(!mem_0_08),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[0]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~6 .extended_lut = "off";
defparam \src_data[0]~6 .lut_mask = 64'hFFCFAA8AF0C0A080;
defparam \src_data[0]~6 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~7 (
	.dataa(!mem_used_018),
	.datab(!mem_0_03),
	.datac(!\src_data[0]~4_combout ),
	.datad(!\src_data[0]~5_combout ),
	.datae(!\src_data[0]~6_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[0]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~7 .extended_lut = "off";
defparam \src_data[0]~7 .lut_mask = 64'h00000E0000000E00;
defparam \src_data[0]~7 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~8 (
	.dataa(!av_readdata_pre_02),
	.datab(!\src_payload~20_combout ),
	.datac(!\src_data[0]~2_combout ),
	.datad(!\src_data[0]~3_combout ),
	.datae(!\src_data[0]~7_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[0]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~8 .extended_lut = "off";
defparam \src_data[0]~8 .lut_mask = 64'h0000E0000000E000;
defparam \src_data[0]~8 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~9 (
	.dataa(!read_latency_shift_reg_02),
	.datab(!mem_used_02),
	.datac(!av_readdata_pre_09),
	.datad(!mem_0_09),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[0]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~9 .extended_lut = "off";
defparam \src_data[0]~9 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[0]~9 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~10 (
	.dataa(!read_latency_shift_reg_03),
	.datab(!mem_used_03),
	.datac(!av_readdata_pre_010),
	.datad(!mem_0_010),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[0]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~10 .extended_lut = "off";
defparam \src_data[0]~10 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[0]~10 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~11 (
	.dataa(!src1_valid1),
	.datab(!src1_valid2),
	.datac(!\src_data[0]~9_combout ),
	.datad(!\src_data[0]~10_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[0]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~11 .extended_lut = "off";
defparam \src_data[0]~11 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[0]~11 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~12 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!av_readdata_pre_011),
	.datad(!mem_0_011),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[0]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~12 .extended_lut = "off";
defparam \src_data[0]~12 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[0]~12 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~13 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_01),
	.datac(!av_readdata_pre_012),
	.datad(!mem_0_012),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[0]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~13 .extended_lut = "off";
defparam \src_data[0]~13 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[0]~13 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~14 (
	.dataa(!read_latency_shift_reg_05),
	.datab(!mem_used_05),
	.datac(!src1_valid7),
	.datad(!av_readdata_pre_013),
	.datae(!mem_0_013),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[0]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~14 .extended_lut = "off";
defparam \src_data[0]~14 .lut_mask = 64'h0040B0F00040B0F0;
defparam \src_data[0]~14 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~15 (
	.dataa(!src1_valid5),
	.datab(!src1_valid6),
	.datac(!\src_data[0]~12_combout ),
	.datad(!\src_data[0]~13_combout ),
	.datae(!\src_data[0]~14_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[0]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~15 .extended_lut = "off";
defparam \src_data[0]~15 .lut_mask = 64'hF5310000F5310000;
defparam \src_data[0]~15 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~16 (
	.dataa(!read_latency_shift_reg_06),
	.datab(!mem_used_06),
	.datac(!av_readdata_pre_014),
	.datad(!mem_0_014),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[0]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~16 .extended_lut = "off";
defparam \src_data[0]~16 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[0]~16 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~17 (
	.dataa(!src1_valid4),
	.datab(!av_readdata_pre_015),
	.datac(!always41),
	.datad(!mem_0_015),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[0]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~17 .extended_lut = "off";
defparam \src_data[0]~17 .lut_mask = 64'h02A202A202A202A2;
defparam \src_data[0]~17 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~18 (
	.dataa(!src1_valid8),
	.datab(!av_readdata_pre_016),
	.datac(!always42),
	.datad(!mem_0_016),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[0]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~18 .extended_lut = "off";
defparam \src_data[0]~18 .lut_mask = 64'h02A202A202A202A2;
defparam \src_data[0]~18 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~19 (
	.dataa(!src1_valid),
	.datab(!\src_data[0]~16_combout ),
	.datac(!\src_data[0]~17_combout ),
	.datad(!\src_data[0]~18_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[0]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~19 .extended_lut = "off";
defparam \src_data[0]~19 .lut_mask = 64'hD000D000D000D000;
defparam \src_data[0]~19 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~23 (
	.dataa(!src1_valid4),
	.datab(!always41),
	.datac(!av_readdata_pre_11),
	.datad(!mem_1_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~23 .extended_lut = "off";
defparam \src_payload~23 .lut_mask = 64'h028A028A028A028A;
defparam \src_payload~23 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~24 (
	.dataa(!read_latency_shift_reg_08),
	.datab(!mem_used_08),
	.datac(!mem_1_02),
	.datad(!av_readdata_pre_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~24 .extended_lut = "off";
defparam \src_payload~24 .lut_mask = 64'h0347034703470347;
defparam \src_payload~24 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~25 (
	.dataa(!mem_used_018),
	.datab(!\src_payload~21_combout ),
	.datac(!av_readdata_pre_13),
	.datad(!mem_1_03),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~25 .extended_lut = "off";
defparam \src_payload~25 .lut_mask = 64'h0357035703570357;
defparam \src_payload~25 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~26 (
	.dataa(!mem_used_016),
	.datab(!\src_payload~22_combout ),
	.datac(!av_readdata_pre_14),
	.datad(!mem_1_04),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~26 .extended_lut = "off";
defparam \src_payload~26 .lut_mask = 64'h0357035703570357;
defparam \src_payload~26 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~27 (
	.dataa(!mem_used_014),
	.datab(!mem_1_01),
	.datac(!\src_payload~24_combout ),
	.datad(!\src_payload~25_combout ),
	.datae(!\src_payload~26_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~27 .extended_lut = "off";
defparam \src_payload~27 .lut_mask = 64'hE0000000E0000000;
defparam \src_payload~27 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~28 (
	.dataa(!src1_valid8),
	.datab(!always42),
	.datac(!av_readdata_pre_15),
	.datad(!mem_1_05),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~28 .extended_lut = "off";
defparam \src_payload~28 .lut_mask = 64'h028A028A028A028A;
defparam \src_payload~28 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~29 (
	.dataa(!src1_valid9),
	.datab(!always4),
	.datac(!\src_payload~28_combout ),
	.datad(!av_readdata_pre_16),
	.datae(!mem_1_06),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~29 .extended_lut = "off";
defparam \src_payload~29 .lut_mask = 64'hF0D07050F0D07050;
defparam \src_payload~29 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~31 (
	.dataa(!src1_valid4),
	.datab(!always41),
	.datac(!av_readdata_pre_21),
	.datad(!mem_2_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~31 .extended_lut = "off";
defparam \src_payload~31 .lut_mask = 64'h028A028A028A028A;
defparam \src_payload~31 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~32 (
	.dataa(!read_latency_shift_reg_08),
	.datab(!mem_used_08),
	.datac(!mem_2_02),
	.datad(!av_readdata_pre_22),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~32 .extended_lut = "off";
defparam \src_payload~32 .lut_mask = 64'h0347034703470347;
defparam \src_payload~32 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~33 (
	.dataa(!mem_used_018),
	.datab(!\src_payload~21_combout ),
	.datac(!av_readdata_pre_23),
	.datad(!mem_2_03),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~33 .extended_lut = "off";
defparam \src_payload~33 .lut_mask = 64'h0357035703570357;
defparam \src_payload~33 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~34 (
	.dataa(!mem_used_016),
	.datab(!\src_payload~22_combout ),
	.datac(!av_readdata_pre_24),
	.datad(!mem_2_04),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~34 .extended_lut = "off";
defparam \src_payload~34 .lut_mask = 64'h0357035703570357;
defparam \src_payload~34 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~35 (
	.dataa(!mem_used_014),
	.datab(!mem_2_01),
	.datac(!\src_payload~32_combout ),
	.datad(!\src_payload~33_combout ),
	.datae(!\src_payload~34_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~35 .extended_lut = "off";
defparam \src_payload~35 .lut_mask = 64'hE0000000E0000000;
defparam \src_payload~35 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~36 (
	.dataa(!src1_valid8),
	.datab(!always42),
	.datac(!av_readdata_pre_25),
	.datad(!mem_2_05),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~36 .extended_lut = "off";
defparam \src_payload~36 .lut_mask = 64'h028A028A028A028A;
defparam \src_payload~36 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~37 (
	.dataa(!src1_valid9),
	.datab(!always4),
	.datac(!\src_payload~36_combout ),
	.datad(!av_readdata_pre_26),
	.datae(!mem_2_06),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~37_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~37 .extended_lut = "off";
defparam \src_payload~37 .lut_mask = 64'hF0D07050F0D07050;
defparam \src_payload~37 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~39 (
	.dataa(!src1_valid4),
	.datab(!always41),
	.datac(!av_readdata_pre_31),
	.datad(!mem_3_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~39 .extended_lut = "off";
defparam \src_payload~39 .lut_mask = 64'h028A028A028A028A;
defparam \src_payload~39 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~40 (
	.dataa(!read_latency_shift_reg_08),
	.datab(!mem_used_08),
	.datac(!mem_3_02),
	.datad(!av_readdata_pre_32),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~40_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~40 .extended_lut = "off";
defparam \src_payload~40 .lut_mask = 64'h0347034703470347;
defparam \src_payload~40 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~41 (
	.dataa(!mem_used_018),
	.datab(!\src_payload~21_combout ),
	.datac(!av_readdata_pre_33),
	.datad(!mem_3_03),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~41_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~41 .extended_lut = "off";
defparam \src_payload~41 .lut_mask = 64'h0357035703570357;
defparam \src_payload~41 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~42 (
	.dataa(!mem_used_014),
	.datab(!mem_3_01),
	.datac(!\src_payload~40_combout ),
	.datad(!\src_payload~41_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~42_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~42 .extended_lut = "off";
defparam \src_payload~42 .lut_mask = 64'hE000E000E000E000;
defparam \src_payload~42 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~43 (
	.dataa(!src1_valid8),
	.datab(!always42),
	.datac(!av_readdata_pre_34),
	.datad(!mem_3_04),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~43_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~43 .extended_lut = "off";
defparam \src_payload~43 .lut_mask = 64'h028A028A028A028A;
defparam \src_payload~43 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~44 (
	.dataa(!src1_valid9),
	.datab(!always4),
	.datac(!\src_payload~43_combout ),
	.datad(!av_readdata_pre_35),
	.datae(!mem_3_05),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~44_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~44 .extended_lut = "off";
defparam \src_payload~44 .lut_mask = 64'hF0D07050F0D07050;
defparam \src_payload~44 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~46 (
	.dataa(!src1_valid4),
	.datab(!always41),
	.datac(!av_readdata_pre_41),
	.datad(!mem_4_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~46_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~46 .extended_lut = "off";
defparam \src_payload~46 .lut_mask = 64'h028A028A028A028A;
defparam \src_payload~46 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~47 (
	.dataa(!read_latency_shift_reg_08),
	.datab(!mem_used_08),
	.datac(!mem_4_02),
	.datad(!av_readdata_pre_42),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~47_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~47 .extended_lut = "off";
defparam \src_payload~47 .lut_mask = 64'h0347034703470347;
defparam \src_payload~47 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~48 (
	.dataa(!mem_used_018),
	.datab(!\src_payload~21_combout ),
	.datac(!av_readdata_pre_43),
	.datad(!mem_4_03),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~48_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~48 .extended_lut = "off";
defparam \src_payload~48 .lut_mask = 64'h0357035703570357;
defparam \src_payload~48 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~49 (
	.dataa(!mem_used_014),
	.datab(!mem_4_01),
	.datac(!\src_payload~47_combout ),
	.datad(!\src_payload~48_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~49_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~49 .extended_lut = "off";
defparam \src_payload~49 .lut_mask = 64'hE000E000E000E000;
defparam \src_payload~49 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~50 (
	.dataa(!src1_valid8),
	.datab(!always42),
	.datac(!av_readdata_pre_44),
	.datad(!mem_4_04),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~50_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~50 .extended_lut = "off";
defparam \src_payload~50 .lut_mask = 64'h028A028A028A028A;
defparam \src_payload~50 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~51 (
	.dataa(!src1_valid9),
	.datab(!always4),
	.datac(!\src_payload~50_combout ),
	.datad(!av_readdata_pre_45),
	.datae(!mem_4_05),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~51_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~51 .extended_lut = "off";
defparam \src_payload~51 .lut_mask = 64'hF0D07050F0D07050;
defparam \src_payload~51 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~53 (
	.dataa(!src1_valid4),
	.datab(!always41),
	.datac(!av_readdata_pre_51),
	.datad(!mem_5_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~53_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~53 .extended_lut = "off";
defparam \src_payload~53 .lut_mask = 64'h028A028A028A028A;
defparam \src_payload~53 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~54 (
	.dataa(!read_latency_shift_reg_08),
	.datab(!mem_used_08),
	.datac(!mem_5_02),
	.datad(!av_readdata_pre_52),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~54_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~54 .extended_lut = "off";
defparam \src_payload~54 .lut_mask = 64'h0347034703470347;
defparam \src_payload~54 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~55 (
	.dataa(!mem_used_018),
	.datab(!\src_payload~21_combout ),
	.datac(!av_readdata_pre_53),
	.datad(!mem_5_03),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~55_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~55 .extended_lut = "off";
defparam \src_payload~55 .lut_mask = 64'h0357035703570357;
defparam \src_payload~55 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~56 (
	.dataa(!mem_used_014),
	.datab(!mem_5_01),
	.datac(!\src_payload~54_combout ),
	.datad(!\src_payload~55_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~56_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~56 .extended_lut = "off";
defparam \src_payload~56 .lut_mask = 64'hE000E000E000E000;
defparam \src_payload~56 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~57 (
	.dataa(!src1_valid8),
	.datab(!always42),
	.datac(!av_readdata_pre_54),
	.datad(!mem_5_04),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~57_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~57 .extended_lut = "off";
defparam \src_payload~57 .lut_mask = 64'h028A028A028A028A;
defparam \src_payload~57 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~58 (
	.dataa(!src1_valid9),
	.datab(!always4),
	.datac(!\src_payload~57_combout ),
	.datad(!av_readdata_pre_55),
	.datae(!mem_5_05),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~58_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~58 .extended_lut = "off";
defparam \src_payload~58 .lut_mask = 64'hF0D07050F0D07050;
defparam \src_payload~58 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~60 (
	.dataa(!src1_valid4),
	.datab(!always41),
	.datac(!av_readdata_pre_61),
	.datad(!mem_6_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~60_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~60 .extended_lut = "off";
defparam \src_payload~60 .lut_mask = 64'h028A028A028A028A;
defparam \src_payload~60 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~61 (
	.dataa(!read_latency_shift_reg_08),
	.datab(!mem_used_08),
	.datac(!mem_6_02),
	.datad(!av_readdata_pre_62),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~61_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~61 .extended_lut = "off";
defparam \src_payload~61 .lut_mask = 64'h0347034703470347;
defparam \src_payload~61 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~62 (
	.dataa(!mem_used_018),
	.datab(!\src_payload~21_combout ),
	.datac(!av_readdata_pre_63),
	.datad(!mem_6_03),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~62_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~62 .extended_lut = "off";
defparam \src_payload~62 .lut_mask = 64'h0357035703570357;
defparam \src_payload~62 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~63 (
	.dataa(!mem_used_014),
	.datab(!mem_6_01),
	.datac(!\src_payload~61_combout ),
	.datad(!\src_payload~62_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~63_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~63 .extended_lut = "off";
defparam \src_payload~63 .lut_mask = 64'hE000E000E000E000;
defparam \src_payload~63 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~64 (
	.dataa(!src1_valid8),
	.datab(!always42),
	.datac(!av_readdata_pre_64),
	.datad(!mem_6_04),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~64_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~64 .extended_lut = "off";
defparam \src_payload~64 .lut_mask = 64'h028A028A028A028A;
defparam \src_payload~64 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~65 (
	.dataa(!src1_valid9),
	.datab(!always4),
	.datac(!\src_payload~64_combout ),
	.datad(!av_readdata_pre_65),
	.datae(!mem_6_05),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~65_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~65 .extended_lut = "off";
defparam \src_payload~65 .lut_mask = 64'hF0D07050F0D07050;
defparam \src_payload~65 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~67 (
	.dataa(!src1_valid4),
	.datab(!always41),
	.datac(!av_readdata_pre_71),
	.datad(!mem_7_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~67_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~67 .extended_lut = "off";
defparam \src_payload~67 .lut_mask = 64'h028A028A028A028A;
defparam \src_payload~67 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~68 (
	.dataa(!src1_valid8),
	.datab(!always42),
	.datac(!av_readdata_pre_72),
	.datad(!mem_7_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~68_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~68 .extended_lut = "off";
defparam \src_payload~68 .lut_mask = 64'h028A028A028A028A;
defparam \src_payload~68 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~69 (
	.dataa(!read_latency_shift_reg_08),
	.datab(!mem_used_08),
	.datac(!mem_7_03),
	.datad(!av_readdata_pre_73),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~69_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~69 .extended_lut = "off";
defparam \src_payload~69 .lut_mask = 64'h0347034703470347;
defparam \src_payload~69 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~70 (
	.dataa(!mem_used_018),
	.datab(!\src_payload~21_combout ),
	.datac(!av_readdata_pre_74),
	.datad(!mem_7_04),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~70_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~70 .extended_lut = "off";
defparam \src_payload~70 .lut_mask = 64'h0357035703570357;
defparam \src_payload~70 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~71 (
	.dataa(!mem_used_014),
	.datab(!mem_7_02),
	.datac(!\src_payload~69_combout ),
	.datad(!\src_payload~70_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~71_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~71 .extended_lut = "off";
defparam \src_payload~71 .lut_mask = 64'hE000E000E000E000;
defparam \src_payload~71 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~73 (
	.dataa(!read_latency_shift_reg_011),
	.datab(!mem_used_014),
	.datac(!mem_8_02),
	.datad(!av_readdata_pre_82),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~73_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~73 .extended_lut = "off";
defparam \src_payload~73 .lut_mask = 64'h0347034703470347;
defparam \src_payload~73 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~74 (
	.dataa(!read_latency_shift_reg_013),
	.datab(!mem_used_018),
	.datac(!mem_8_01),
	.datad(!av_readdata_pre_81),
	.datae(!\src_payload~73_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~74_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~74 .extended_lut = "off";
defparam \src_payload~74 .lut_mask = 64'hFCB80000FCB80000;
defparam \src_payload~74 .shared_arith = "off";

cyclonev_lcell_comb \src_data[105]~21 (
	.dataa(!empty5),
	.datab(!empty6),
	.datac(!mem_105_011),
	.datad(!mem_105_012),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[105]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[105]~21 .extended_lut = "off";
defparam \src_data[105]~21 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[105]~21 .shared_arith = "off";

cyclonev_lcell_comb \src_data[105]~22 (
	.dataa(!empty),
	.datab(!empty4),
	.datac(!mem_105_013),
	.datad(!mem_105_014),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[105]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[105]~22 .extended_lut = "off";
defparam \src_data[105]~22 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[105]~22 .shared_arith = "off";

cyclonev_lcell_comb \src_data[105]~23 (
	.dataa(!empty3),
	.datab(!empty2),
	.datac(!mem_105_015),
	.datad(!mem_105_016),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[105]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[105]~23 .extended_lut = "off";
defparam \src_data[105]~23 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[105]~23 .shared_arith = "off";

cyclonev_lcell_comb \src_data[105]~24 (
	.dataa(!src1_valid1),
	.datab(!mem_105_06),
	.datac(!\src_data[105]~21_combout ),
	.datad(!\src_data[105]~22_combout ),
	.datae(!\src_data[105]~23_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[105]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[105]~24 .extended_lut = "off";
defparam \src_data[105]~24 .lut_mask = 64'hD0000000D0000000;
defparam \src_data[105]~24 .shared_arith = "off";

cyclonev_lcell_comb \src_data[105]~25 (
	.dataa(!src1_valid2),
	.datab(!src1_valid3),
	.datac(!src1_valid4),
	.datad(!mem_105_07),
	.datae(!mem_105_04),
	.dataf(!mem_105_08),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[105]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[105]~25 .extended_lut = "off";
defparam \src_data[105]~25 .lut_mask = 64'hFF5533110F050301;
defparam \src_data[105]~25 .shared_arith = "off";

cyclonev_lcell_comb \src_data[105]~26 (
	.dataa(!src1_valid5),
	.datab(!src1_valid6),
	.datac(!src1_valid7),
	.datad(!mem_105_09),
	.datae(!mem_105_05),
	.dataf(!mem_105_02),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[105]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[105]~26 .extended_lut = "off";
defparam \src_data[105]~26 .lut_mask = 64'hFF5533110F050301;
defparam \src_data[105]~26 .shared_arith = "off";

cyclonev_lcell_comb \src_data[105]~27 (
	.dataa(!src1_valid8),
	.datab(!src1_valid9),
	.datac(!src1_valid),
	.datad(!mem_105_03),
	.datae(!mem_105_0),
	.dataf(!mem_105_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[105]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[105]~27 .extended_lut = "off";
defparam \src_data[105]~27 .lut_mask = 64'hFF5533110F050301;
defparam \src_data[105]~27 .shared_arith = "off";

cyclonev_lcell_comb \src_data[106]~28 (
	.dataa(!empty5),
	.datab(!empty6),
	.datac(!mem_106_011),
	.datad(!mem_106_012),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[106]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[106]~28 .extended_lut = "off";
defparam \src_data[106]~28 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[106]~28 .shared_arith = "off";

cyclonev_lcell_comb \src_data[106]~29 (
	.dataa(!empty),
	.datab(!empty4),
	.datac(!mem_106_013),
	.datad(!mem_106_014),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[106]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[106]~29 .extended_lut = "off";
defparam \src_data[106]~29 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[106]~29 .shared_arith = "off";

cyclonev_lcell_comb \src_data[106]~30 (
	.dataa(!empty3),
	.datab(!empty2),
	.datac(!mem_106_015),
	.datad(!mem_106_016),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[106]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[106]~30 .extended_lut = "off";
defparam \src_data[106]~30 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[106]~30 .shared_arith = "off";

cyclonev_lcell_comb \src_data[106]~31 (
	.dataa(!src1_valid1),
	.datab(!mem_106_06),
	.datac(!\src_data[106]~28_combout ),
	.datad(!\src_data[106]~29_combout ),
	.datae(!\src_data[106]~30_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[106]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[106]~31 .extended_lut = "off";
defparam \src_data[106]~31 .lut_mask = 64'hD0000000D0000000;
defparam \src_data[106]~31 .shared_arith = "off";

cyclonev_lcell_comb \src_data[106]~32 (
	.dataa(!src1_valid2),
	.datab(!src1_valid3),
	.datac(!src1_valid4),
	.datad(!mem_106_07),
	.datae(!mem_106_04),
	.dataf(!mem_106_08),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[106]~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[106]~32 .extended_lut = "off";
defparam \src_data[106]~32 .lut_mask = 64'hFF5533110F050301;
defparam \src_data[106]~32 .shared_arith = "off";

cyclonev_lcell_comb \src_data[106]~33 (
	.dataa(!src1_valid5),
	.datab(!src1_valid6),
	.datac(!src1_valid7),
	.datad(!mem_106_09),
	.datae(!mem_106_05),
	.dataf(!mem_106_02),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[106]~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[106]~33 .extended_lut = "off";
defparam \src_data[106]~33 .lut_mask = 64'hFF5533110F050301;
defparam \src_data[106]~33 .shared_arith = "off";

cyclonev_lcell_comb \src_data[106]~34 (
	.dataa(!src1_valid8),
	.datab(!src1_valid9),
	.datac(!src1_valid),
	.datad(!mem_106_03),
	.datae(!mem_106_0),
	.dataf(!mem_106_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[106]~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[106]~34 .extended_lut = "off";
defparam \src_data[106]~34 .lut_mask = 64'hFF5533110F050301;
defparam \src_data[106]~34 .shared_arith = "off";

cyclonev_lcell_comb \src_data[107]~35 (
	.dataa(!empty5),
	.datab(!empty6),
	.datac(!mem_107_011),
	.datad(!mem_107_012),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[107]~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[107]~35 .extended_lut = "off";
defparam \src_data[107]~35 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[107]~35 .shared_arith = "off";

cyclonev_lcell_comb \src_data[107]~36 (
	.dataa(!empty),
	.datab(!empty4),
	.datac(!mem_107_013),
	.datad(!mem_107_014),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[107]~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[107]~36 .extended_lut = "off";
defparam \src_data[107]~36 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[107]~36 .shared_arith = "off";

cyclonev_lcell_comb \src_data[107]~37 (
	.dataa(!empty3),
	.datab(!empty2),
	.datac(!mem_107_015),
	.datad(!mem_107_016),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[107]~37_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[107]~37 .extended_lut = "off";
defparam \src_data[107]~37 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[107]~37 .shared_arith = "off";

cyclonev_lcell_comb \src_data[107]~38 (
	.dataa(!src1_valid1),
	.datab(!mem_107_06),
	.datac(!\src_data[107]~35_combout ),
	.datad(!\src_data[107]~36_combout ),
	.datae(!\src_data[107]~37_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[107]~38_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[107]~38 .extended_lut = "off";
defparam \src_data[107]~38 .lut_mask = 64'hD0000000D0000000;
defparam \src_data[107]~38 .shared_arith = "off";

cyclonev_lcell_comb \src_data[107]~39 (
	.dataa(!src1_valid2),
	.datab(!src1_valid3),
	.datac(!src1_valid4),
	.datad(!mem_107_07),
	.datae(!mem_107_04),
	.dataf(!mem_107_08),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[107]~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[107]~39 .extended_lut = "off";
defparam \src_data[107]~39 .lut_mask = 64'hFF5533110F050301;
defparam \src_data[107]~39 .shared_arith = "off";

cyclonev_lcell_comb \src_data[107]~40 (
	.dataa(!src1_valid5),
	.datab(!src1_valid6),
	.datac(!src1_valid7),
	.datad(!mem_107_09),
	.datae(!mem_107_05),
	.dataf(!mem_107_02),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[107]~40_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[107]~40 .extended_lut = "off";
defparam \src_data[107]~40 .lut_mask = 64'hFF5533110F050301;
defparam \src_data[107]~40 .shared_arith = "off";

cyclonev_lcell_comb \src_data[107]~41 (
	.dataa(!src1_valid8),
	.datab(!src1_valid9),
	.datac(!src1_valid),
	.datad(!mem_107_03),
	.datae(!mem_107_0),
	.dataf(!mem_107_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[107]~41_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[107]~41 .extended_lut = "off";
defparam \src_data[107]~41 .lut_mask = 64'hFF5533110F050301;
defparam \src_data[107]~41 .shared_arith = "off";

cyclonev_lcell_comb \src_data[108]~42 (
	.dataa(!empty5),
	.datab(!empty6),
	.datac(!mem_108_011),
	.datad(!mem_108_012),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[108]~42_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[108]~42 .extended_lut = "off";
defparam \src_data[108]~42 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[108]~42 .shared_arith = "off";

cyclonev_lcell_comb \src_data[108]~43 (
	.dataa(!empty),
	.datab(!empty4),
	.datac(!mem_108_013),
	.datad(!mem_108_014),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[108]~43_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[108]~43 .extended_lut = "off";
defparam \src_data[108]~43 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[108]~43 .shared_arith = "off";

cyclonev_lcell_comb \src_data[108]~44 (
	.dataa(!empty3),
	.datab(!empty2),
	.datac(!mem_108_015),
	.datad(!mem_108_016),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[108]~44_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[108]~44 .extended_lut = "off";
defparam \src_data[108]~44 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[108]~44 .shared_arith = "off";

cyclonev_lcell_comb \src_data[108]~45 (
	.dataa(!src1_valid1),
	.datab(!mem_108_06),
	.datac(!\src_data[108]~42_combout ),
	.datad(!\src_data[108]~43_combout ),
	.datae(!\src_data[108]~44_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[108]~45_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[108]~45 .extended_lut = "off";
defparam \src_data[108]~45 .lut_mask = 64'hD0000000D0000000;
defparam \src_data[108]~45 .shared_arith = "off";

cyclonev_lcell_comb \src_data[108]~46 (
	.dataa(!src1_valid2),
	.datab(!src1_valid3),
	.datac(!src1_valid4),
	.datad(!mem_108_07),
	.datae(!mem_108_04),
	.dataf(!mem_108_08),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[108]~46_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[108]~46 .extended_lut = "off";
defparam \src_data[108]~46 .lut_mask = 64'hFF5533110F050301;
defparam \src_data[108]~46 .shared_arith = "off";

cyclonev_lcell_comb \src_data[108]~47 (
	.dataa(!src1_valid5),
	.datab(!src1_valid6),
	.datac(!src1_valid7),
	.datad(!mem_108_09),
	.datae(!mem_108_05),
	.dataf(!mem_108_02),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[108]~47_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[108]~47 .extended_lut = "off";
defparam \src_data[108]~47 .lut_mask = 64'hFF5533110F050301;
defparam \src_data[108]~47 .shared_arith = "off";

cyclonev_lcell_comb \src_data[108]~48 (
	.dataa(!src1_valid8),
	.datab(!src1_valid9),
	.datac(!src1_valid),
	.datad(!mem_108_03),
	.datae(!mem_108_0),
	.dataf(!mem_108_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[108]~48_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[108]~48 .extended_lut = "off";
defparam \src_data[108]~48 .lut_mask = 64'hFF5533110F050301;
defparam \src_data[108]~48 .shared_arith = "off";

cyclonev_lcell_comb \src_data[109]~49 (
	.dataa(!empty5),
	.datab(!empty6),
	.datac(!mem_109_011),
	.datad(!mem_109_012),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[109]~49_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[109]~49 .extended_lut = "off";
defparam \src_data[109]~49 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[109]~49 .shared_arith = "off";

cyclonev_lcell_comb \src_data[109]~50 (
	.dataa(!empty),
	.datab(!empty4),
	.datac(!mem_109_013),
	.datad(!mem_109_014),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[109]~50_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[109]~50 .extended_lut = "off";
defparam \src_data[109]~50 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[109]~50 .shared_arith = "off";

cyclonev_lcell_comb \src_data[109]~51 (
	.dataa(!empty3),
	.datab(!empty2),
	.datac(!mem_109_015),
	.datad(!mem_109_016),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[109]~51_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[109]~51 .extended_lut = "off";
defparam \src_data[109]~51 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[109]~51 .shared_arith = "off";

cyclonev_lcell_comb \src_data[109]~52 (
	.dataa(!src1_valid1),
	.datab(!mem_109_06),
	.datac(!\src_data[109]~49_combout ),
	.datad(!\src_data[109]~50_combout ),
	.datae(!\src_data[109]~51_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[109]~52_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[109]~52 .extended_lut = "off";
defparam \src_data[109]~52 .lut_mask = 64'hD0000000D0000000;
defparam \src_data[109]~52 .shared_arith = "off";

cyclonev_lcell_comb \src_data[109]~53 (
	.dataa(!src1_valid2),
	.datab(!src1_valid3),
	.datac(!src1_valid4),
	.datad(!mem_109_07),
	.datae(!mem_109_04),
	.dataf(!mem_109_08),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[109]~53_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[109]~53 .extended_lut = "off";
defparam \src_data[109]~53 .lut_mask = 64'hFF5533110F050301;
defparam \src_data[109]~53 .shared_arith = "off";

cyclonev_lcell_comb \src_data[109]~54 (
	.dataa(!src1_valid5),
	.datab(!src1_valid6),
	.datac(!src1_valid7),
	.datad(!mem_109_09),
	.datae(!mem_109_05),
	.dataf(!mem_109_02),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[109]~54_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[109]~54 .extended_lut = "off";
defparam \src_data[109]~54 .lut_mask = 64'hFF5533110F050301;
defparam \src_data[109]~54 .shared_arith = "off";

cyclonev_lcell_comb \src_data[109]~55 (
	.dataa(!src1_valid8),
	.datab(!src1_valid9),
	.datac(!src1_valid),
	.datad(!mem_109_03),
	.datae(!mem_109_0),
	.dataf(!mem_109_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[109]~55_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[109]~55 .extended_lut = "off";
defparam \src_data[109]~55 .lut_mask = 64'hFF5533110F050301;
defparam \src_data[109]~55 .shared_arith = "off";

cyclonev_lcell_comb \src_data[110]~56 (
	.dataa(!empty5),
	.datab(!empty6),
	.datac(!mem_110_011),
	.datad(!mem_110_012),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[110]~56_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[110]~56 .extended_lut = "off";
defparam \src_data[110]~56 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[110]~56 .shared_arith = "off";

cyclonev_lcell_comb \src_data[110]~57 (
	.dataa(!empty),
	.datab(!empty4),
	.datac(!mem_110_013),
	.datad(!mem_110_014),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[110]~57_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[110]~57 .extended_lut = "off";
defparam \src_data[110]~57 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[110]~57 .shared_arith = "off";

cyclonev_lcell_comb \src_data[110]~58 (
	.dataa(!empty3),
	.datab(!empty2),
	.datac(!mem_110_015),
	.datad(!mem_110_016),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[110]~58_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[110]~58 .extended_lut = "off";
defparam \src_data[110]~58 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[110]~58 .shared_arith = "off";

cyclonev_lcell_comb \src_data[110]~59 (
	.dataa(!src1_valid1),
	.datab(!mem_110_06),
	.datac(!\src_data[110]~56_combout ),
	.datad(!\src_data[110]~57_combout ),
	.datae(!\src_data[110]~58_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[110]~59_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[110]~59 .extended_lut = "off";
defparam \src_data[110]~59 .lut_mask = 64'hD0000000D0000000;
defparam \src_data[110]~59 .shared_arith = "off";

cyclonev_lcell_comb \src_data[110]~60 (
	.dataa(!src1_valid2),
	.datab(!src1_valid3),
	.datac(!src1_valid4),
	.datad(!mem_110_07),
	.datae(!mem_110_04),
	.dataf(!mem_110_08),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[110]~60_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[110]~60 .extended_lut = "off";
defparam \src_data[110]~60 .lut_mask = 64'hFF5533110F050301;
defparam \src_data[110]~60 .shared_arith = "off";

cyclonev_lcell_comb \src_data[110]~61 (
	.dataa(!src1_valid5),
	.datab(!src1_valid6),
	.datac(!src1_valid7),
	.datad(!mem_110_09),
	.datae(!mem_110_05),
	.dataf(!mem_110_02),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[110]~61_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[110]~61 .extended_lut = "off";
defparam \src_data[110]~61 .lut_mask = 64'hFF5533110F050301;
defparam \src_data[110]~61 .shared_arith = "off";

cyclonev_lcell_comb \src_data[110]~62 (
	.dataa(!src1_valid8),
	.datab(!src1_valid9),
	.datac(!src1_valid),
	.datad(!mem_110_03),
	.datae(!mem_110_0),
	.dataf(!mem_110_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[110]~62_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[110]~62 .extended_lut = "off";
defparam \src_data[110]~62 .lut_mask = 64'hFF5533110F050301;
defparam \src_data[110]~62 .shared_arith = "off";

cyclonev_lcell_comb \src_data[111]~63 (
	.dataa(!empty5),
	.datab(!empty6),
	.datac(!mem_111_011),
	.datad(!mem_111_012),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[111]~63_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[111]~63 .extended_lut = "off";
defparam \src_data[111]~63 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[111]~63 .shared_arith = "off";

cyclonev_lcell_comb \src_data[111]~64 (
	.dataa(!empty),
	.datab(!empty4),
	.datac(!mem_111_013),
	.datad(!mem_111_014),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[111]~64_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[111]~64 .extended_lut = "off";
defparam \src_data[111]~64 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[111]~64 .shared_arith = "off";

cyclonev_lcell_comb \src_data[111]~65 (
	.dataa(!empty3),
	.datab(!empty2),
	.datac(!mem_111_015),
	.datad(!mem_111_016),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[111]~65_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[111]~65 .extended_lut = "off";
defparam \src_data[111]~65 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[111]~65 .shared_arith = "off";

cyclonev_lcell_comb \src_data[111]~66 (
	.dataa(!src1_valid1),
	.datab(!mem_111_06),
	.datac(!\src_data[111]~63_combout ),
	.datad(!\src_data[111]~64_combout ),
	.datae(!\src_data[111]~65_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[111]~66_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[111]~66 .extended_lut = "off";
defparam \src_data[111]~66 .lut_mask = 64'hD0000000D0000000;
defparam \src_data[111]~66 .shared_arith = "off";

cyclonev_lcell_comb \src_data[111]~67 (
	.dataa(!src1_valid2),
	.datab(!src1_valid3),
	.datac(!src1_valid4),
	.datad(!mem_111_07),
	.datae(!mem_111_04),
	.dataf(!mem_111_08),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[111]~67_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[111]~67 .extended_lut = "off";
defparam \src_data[111]~67 .lut_mask = 64'hFF5533110F050301;
defparam \src_data[111]~67 .shared_arith = "off";

cyclonev_lcell_comb \src_data[111]~68 (
	.dataa(!src1_valid5),
	.datab(!src1_valid6),
	.datac(!src1_valid7),
	.datad(!mem_111_09),
	.datae(!mem_111_05),
	.dataf(!mem_111_02),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[111]~68_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[111]~68 .extended_lut = "off";
defparam \src_data[111]~68 .lut_mask = 64'hFF5533110F050301;
defparam \src_data[111]~68 .shared_arith = "off";

cyclonev_lcell_comb \src_data[111]~69 (
	.dataa(!src1_valid8),
	.datab(!src1_valid9),
	.datac(!src1_valid),
	.datad(!mem_111_03),
	.datae(!mem_111_0),
	.dataf(!mem_111_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[111]~69_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[111]~69 .extended_lut = "off";
defparam \src_data[111]~69 .lut_mask = 64'hFF5533110F050301;
defparam \src_data[111]~69 .shared_arith = "off";

cyclonev_lcell_comb \src_data[112]~70 (
	.dataa(!empty5),
	.datab(!empty6),
	.datac(!mem_112_011),
	.datad(!mem_112_012),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[112]~70_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[112]~70 .extended_lut = "off";
defparam \src_data[112]~70 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[112]~70 .shared_arith = "off";

cyclonev_lcell_comb \src_data[112]~71 (
	.dataa(!empty),
	.datab(!empty4),
	.datac(!mem_112_013),
	.datad(!mem_112_014),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[112]~71_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[112]~71 .extended_lut = "off";
defparam \src_data[112]~71 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[112]~71 .shared_arith = "off";

cyclonev_lcell_comb \src_data[112]~72 (
	.dataa(!empty3),
	.datab(!empty2),
	.datac(!mem_112_015),
	.datad(!mem_112_016),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[112]~72_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[112]~72 .extended_lut = "off";
defparam \src_data[112]~72 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[112]~72 .shared_arith = "off";

cyclonev_lcell_comb \src_data[112]~73 (
	.dataa(!src1_valid1),
	.datab(!mem_112_06),
	.datac(!\src_data[112]~70_combout ),
	.datad(!\src_data[112]~71_combout ),
	.datae(!\src_data[112]~72_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[112]~73_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[112]~73 .extended_lut = "off";
defparam \src_data[112]~73 .lut_mask = 64'hD0000000D0000000;
defparam \src_data[112]~73 .shared_arith = "off";

cyclonev_lcell_comb \src_data[112]~74 (
	.dataa(!src1_valid2),
	.datab(!src1_valid3),
	.datac(!src1_valid4),
	.datad(!mem_112_07),
	.datae(!mem_112_04),
	.dataf(!mem_112_08),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[112]~74_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[112]~74 .extended_lut = "off";
defparam \src_data[112]~74 .lut_mask = 64'hFF5533110F050301;
defparam \src_data[112]~74 .shared_arith = "off";

cyclonev_lcell_comb \src_data[112]~75 (
	.dataa(!src1_valid5),
	.datab(!src1_valid6),
	.datac(!src1_valid7),
	.datad(!mem_112_09),
	.datae(!mem_112_05),
	.dataf(!mem_112_02),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[112]~75_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[112]~75 .extended_lut = "off";
defparam \src_data[112]~75 .lut_mask = 64'hFF5533110F050301;
defparam \src_data[112]~75 .shared_arith = "off";

cyclonev_lcell_comb \src_data[112]~76 (
	.dataa(!src1_valid8),
	.datab(!src1_valid9),
	.datac(!src1_valid),
	.datad(!mem_112_03),
	.datae(!mem_112_0),
	.dataf(!mem_112_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[112]~76_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[112]~76 .extended_lut = "off";
defparam \src_data[112]~76 .lut_mask = 64'hFF5533110F050301;
defparam \src_data[112]~76 .shared_arith = "off";

cyclonev_lcell_comb \src_data[113]~77 (
	.dataa(!empty5),
	.datab(!empty6),
	.datac(!mem_113_011),
	.datad(!mem_113_012),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[113]~77_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[113]~77 .extended_lut = "off";
defparam \src_data[113]~77 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[113]~77 .shared_arith = "off";

cyclonev_lcell_comb \src_data[113]~78 (
	.dataa(!empty),
	.datab(!empty4),
	.datac(!mem_113_013),
	.datad(!mem_113_014),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[113]~78_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[113]~78 .extended_lut = "off";
defparam \src_data[113]~78 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[113]~78 .shared_arith = "off";

cyclonev_lcell_comb \src_data[113]~79 (
	.dataa(!empty3),
	.datab(!empty2),
	.datac(!mem_113_015),
	.datad(!mem_113_016),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[113]~79_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[113]~79 .extended_lut = "off";
defparam \src_data[113]~79 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[113]~79 .shared_arith = "off";

cyclonev_lcell_comb \src_data[113]~80 (
	.dataa(!src1_valid1),
	.datab(!mem_113_06),
	.datac(!\src_data[113]~77_combout ),
	.datad(!\src_data[113]~78_combout ),
	.datae(!\src_data[113]~79_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[113]~80_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[113]~80 .extended_lut = "off";
defparam \src_data[113]~80 .lut_mask = 64'hD0000000D0000000;
defparam \src_data[113]~80 .shared_arith = "off";

cyclonev_lcell_comb \src_data[113]~81 (
	.dataa(!src1_valid2),
	.datab(!src1_valid3),
	.datac(!src1_valid4),
	.datad(!mem_113_07),
	.datae(!mem_113_04),
	.dataf(!mem_113_08),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[113]~81_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[113]~81 .extended_lut = "off";
defparam \src_data[113]~81 .lut_mask = 64'hFF5533110F050301;
defparam \src_data[113]~81 .shared_arith = "off";

cyclonev_lcell_comb \src_data[113]~82 (
	.dataa(!src1_valid5),
	.datab(!src1_valid6),
	.datac(!src1_valid7),
	.datad(!mem_113_09),
	.datae(!mem_113_05),
	.dataf(!mem_113_02),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[113]~82_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[113]~82 .extended_lut = "off";
defparam \src_data[113]~82 .lut_mask = 64'hFF5533110F050301;
defparam \src_data[113]~82 .shared_arith = "off";

cyclonev_lcell_comb \src_data[113]~83 (
	.dataa(!src1_valid8),
	.datab(!src1_valid9),
	.datac(!src1_valid),
	.datad(!mem_113_03),
	.datae(!mem_113_0),
	.dataf(!mem_113_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[113]~83_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[113]~83 .extended_lut = "off";
defparam \src_data[113]~83 .lut_mask = 64'hFF5533110F050301;
defparam \src_data[113]~83 .shared_arith = "off";

cyclonev_lcell_comb \src_data[114]~84 (
	.dataa(!empty5),
	.datab(!empty6),
	.datac(!mem_114_011),
	.datad(!mem_114_012),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[114]~84_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[114]~84 .extended_lut = "off";
defparam \src_data[114]~84 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[114]~84 .shared_arith = "off";

cyclonev_lcell_comb \src_data[114]~85 (
	.dataa(!empty),
	.datab(!empty4),
	.datac(!mem_114_013),
	.datad(!mem_114_014),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[114]~85_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[114]~85 .extended_lut = "off";
defparam \src_data[114]~85 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[114]~85 .shared_arith = "off";

cyclonev_lcell_comb \src_data[114]~86 (
	.dataa(!empty3),
	.datab(!empty2),
	.datac(!mem_114_015),
	.datad(!mem_114_016),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[114]~86_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[114]~86 .extended_lut = "off";
defparam \src_data[114]~86 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[114]~86 .shared_arith = "off";

cyclonev_lcell_comb \src_data[114]~87 (
	.dataa(!src1_valid1),
	.datab(!mem_114_06),
	.datac(!\src_data[114]~84_combout ),
	.datad(!\src_data[114]~85_combout ),
	.datae(!\src_data[114]~86_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[114]~87_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[114]~87 .extended_lut = "off";
defparam \src_data[114]~87 .lut_mask = 64'hD0000000D0000000;
defparam \src_data[114]~87 .shared_arith = "off";

cyclonev_lcell_comb \src_data[114]~88 (
	.dataa(!src1_valid2),
	.datab(!src1_valid3),
	.datac(!src1_valid4),
	.datad(!mem_114_07),
	.datae(!mem_114_04),
	.dataf(!mem_114_08),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[114]~88_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[114]~88 .extended_lut = "off";
defparam \src_data[114]~88 .lut_mask = 64'hFF5533110F050301;
defparam \src_data[114]~88 .shared_arith = "off";

cyclonev_lcell_comb \src_data[114]~89 (
	.dataa(!src1_valid5),
	.datab(!src1_valid6),
	.datac(!src1_valid7),
	.datad(!mem_114_09),
	.datae(!mem_114_05),
	.dataf(!mem_114_02),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[114]~89_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[114]~89 .extended_lut = "off";
defparam \src_data[114]~89 .lut_mask = 64'hFF5533110F050301;
defparam \src_data[114]~89 .shared_arith = "off";

cyclonev_lcell_comb \src_data[114]~90 (
	.dataa(!src1_valid8),
	.datab(!src1_valid9),
	.datac(!src1_valid),
	.datad(!mem_114_03),
	.datae(!mem_114_0),
	.dataf(!mem_114_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[114]~90_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[114]~90 .extended_lut = "off";
defparam \src_data[114]~90 .lut_mask = 64'hFF5533110F050301;
defparam \src_data[114]~90 .shared_arith = "off";

cyclonev_lcell_comb \src_data[115]~91 (
	.dataa(!empty5),
	.datab(!empty6),
	.datac(!mem_115_011),
	.datad(!mem_115_012),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[115]~91_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[115]~91 .extended_lut = "off";
defparam \src_data[115]~91 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[115]~91 .shared_arith = "off";

cyclonev_lcell_comb \src_data[115]~92 (
	.dataa(!empty),
	.datab(!empty4),
	.datac(!mem_115_013),
	.datad(!mem_115_014),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[115]~92_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[115]~92 .extended_lut = "off";
defparam \src_data[115]~92 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[115]~92 .shared_arith = "off";

cyclonev_lcell_comb \src_data[115]~93 (
	.dataa(!empty3),
	.datab(!empty2),
	.datac(!mem_115_015),
	.datad(!mem_115_016),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[115]~93_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[115]~93 .extended_lut = "off";
defparam \src_data[115]~93 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[115]~93 .shared_arith = "off";

cyclonev_lcell_comb \src_data[115]~94 (
	.dataa(!src1_valid1),
	.datab(!mem_115_06),
	.datac(!\src_data[115]~91_combout ),
	.datad(!\src_data[115]~92_combout ),
	.datae(!\src_data[115]~93_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[115]~94_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[115]~94 .extended_lut = "off";
defparam \src_data[115]~94 .lut_mask = 64'hD0000000D0000000;
defparam \src_data[115]~94 .shared_arith = "off";

cyclonev_lcell_comb \src_data[115]~95 (
	.dataa(!src1_valid2),
	.datab(!src1_valid3),
	.datac(!src1_valid4),
	.datad(!mem_115_07),
	.datae(!mem_115_04),
	.dataf(!mem_115_08),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[115]~95_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[115]~95 .extended_lut = "off";
defparam \src_data[115]~95 .lut_mask = 64'hFF5533110F050301;
defparam \src_data[115]~95 .shared_arith = "off";

cyclonev_lcell_comb \src_data[115]~96 (
	.dataa(!src1_valid5),
	.datab(!src1_valid6),
	.datac(!src1_valid7),
	.datad(!mem_115_09),
	.datae(!mem_115_05),
	.dataf(!mem_115_02),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[115]~96_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[115]~96 .extended_lut = "off";
defparam \src_data[115]~96 .lut_mask = 64'hFF5533110F050301;
defparam \src_data[115]~96 .shared_arith = "off";

cyclonev_lcell_comb \src_data[115]~97 (
	.dataa(!src1_valid8),
	.datab(!src1_valid9),
	.datac(!src1_valid),
	.datad(!mem_115_03),
	.datae(!mem_115_0),
	.dataf(!mem_115_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[115]~97_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[115]~97 .extended_lut = "off";
defparam \src_data[115]~97 .lut_mask = 64'hFF5533110F050301;
defparam \src_data[115]~97 .shared_arith = "off";

cyclonev_lcell_comb \src_data[116]~98 (
	.dataa(!empty5),
	.datab(!empty6),
	.datac(!mem_116_011),
	.datad(!mem_116_012),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[116]~98_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[116]~98 .extended_lut = "off";
defparam \src_data[116]~98 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[116]~98 .shared_arith = "off";

cyclonev_lcell_comb \src_data[116]~99 (
	.dataa(!empty),
	.datab(!empty4),
	.datac(!mem_116_013),
	.datad(!mem_116_014),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[116]~99_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[116]~99 .extended_lut = "off";
defparam \src_data[116]~99 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[116]~99 .shared_arith = "off";

cyclonev_lcell_comb \src_data[116]~100 (
	.dataa(!empty3),
	.datab(!empty2),
	.datac(!mem_116_015),
	.datad(!mem_116_016),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[116]~100_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[116]~100 .extended_lut = "off";
defparam \src_data[116]~100 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[116]~100 .shared_arith = "off";

cyclonev_lcell_comb \src_data[116]~101 (
	.dataa(!src1_valid1),
	.datab(!mem_116_06),
	.datac(!\src_data[116]~98_combout ),
	.datad(!\src_data[116]~99_combout ),
	.datae(!\src_data[116]~100_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[116]~101_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[116]~101 .extended_lut = "off";
defparam \src_data[116]~101 .lut_mask = 64'hD0000000D0000000;
defparam \src_data[116]~101 .shared_arith = "off";

cyclonev_lcell_comb \src_data[116]~102 (
	.dataa(!src1_valid2),
	.datab(!src1_valid3),
	.datac(!src1_valid4),
	.datad(!mem_116_07),
	.datae(!mem_116_04),
	.dataf(!mem_116_08),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[116]~102_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[116]~102 .extended_lut = "off";
defparam \src_data[116]~102 .lut_mask = 64'hFF5533110F050301;
defparam \src_data[116]~102 .shared_arith = "off";

cyclonev_lcell_comb \src_data[116]~103 (
	.dataa(!src1_valid5),
	.datab(!src1_valid6),
	.datac(!src1_valid7),
	.datad(!mem_116_09),
	.datae(!mem_116_05),
	.dataf(!mem_116_02),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[116]~103_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[116]~103 .extended_lut = "off";
defparam \src_data[116]~103 .lut_mask = 64'hFF5533110F050301;
defparam \src_data[116]~103 .shared_arith = "off";

cyclonev_lcell_comb \src_data[116]~104 (
	.dataa(!src1_valid8),
	.datab(!src1_valid9),
	.datac(!src1_valid),
	.datad(!mem_116_03),
	.datae(!mem_116_0),
	.dataf(!mem_116_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[116]~104_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[116]~104 .extended_lut = "off";
defparam \src_data[116]~104 .lut_mask = 64'hFF5533110F050301;
defparam \src_data[116]~104 .shared_arith = "off";

endmodule

module spw_babasu_spw_babasu_pll_0 (
	outclk_wire_0,
	locked,
	clk_clk,
	reset_reset_n)/* synthesis synthesis_greybox=0 */;
output 	outclk_wire_0;
output 	locked;
input 	clk_clk;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



spw_babasu_altera_pll_1 altera_pll_i(
	.outclk({outclk_wire_0}),
	.locked(locked),
	.refclk(clk_clk),
	.rst(reset_reset_n));

endmodule

module spw_babasu_altera_pll_1 (
	outclk,
	locked,
	refclk,
	rst)/* synthesis synthesis_greybox=0 */;
output 	[0:0] outclk;
output 	locked;
input 	refclk;
input 	rst;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fboutclk_wire[0] ;


generic_pll \general[0].gpll (
	.refclk(refclk),
	.fbclk(\fboutclk_wire[0] ),
	.rst(!rst),
	.writerefclkdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.writeoutclkdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.writephaseshiftdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.writedutycycledata(64'b0000000000000000000000000000000000000000000000000000000000000000),
	.outclk(outclk[0]),
	.fboutclk(\fboutclk_wire[0] ),
	.locked(locked),
	.readrefclkdata(),
	.readoutclkdata(),
	.readphaseshiftdata(),
	.readdutycycledata());
defparam \general[0].gpll .clock_name_global = "false";
defparam \general[0].gpll .duty_cycle = 50;
defparam \general[0].gpll .fractional_vco_multiplier = "false";
defparam \general[0].gpll .output_clock_frequency = "200.0 mhz";
defparam \general[0].gpll .phase_shift = "0 ps";
defparam \general[0].gpll .reference_clock_frequency = "50.0 mhz";
defparam \general[0].gpll .simulation_type = "timing";

endmodule

module spw_babasu_spw_babasu_RX_EMPTY (
	altera_reset_synchronizer_int_chain_out,
	readdata_0,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	clk_clk,
	rx_empty_external_connection_export)/* synthesis synthesis_greybox=0 */;
input 	altera_reset_synchronizer_int_chain_out;
output 	readdata_0;
input 	int_nxt_addr_reg_dly_3;
input 	int_nxt_addr_reg_dly_2;
input 	clk_clk;
input 	rx_empty_external_connection_export;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_mux_out~combout ;


dffeas \readdata[0] (
	.clk(clk_clk),
	.d(\read_mux_out~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

cyclonev_lcell_comb read_mux_out(
	.dataa(!rx_empty_external_connection_export),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam read_mux_out.extended_lut = "off";
defparam read_mux_out.lut_mask = 64'h4040404040404040;
defparam read_mux_out.shared_arith = "off";

endmodule

module spw_babasu_spw_babasu_RX_EMPTY_1 (
	altera_reset_synchronizer_int_chain_out,
	readdata_0,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	clk_clk,
	tick_out_external_connection_export)/* synthesis synthesis_greybox=0 */;
input 	altera_reset_synchronizer_int_chain_out;
output 	readdata_0;
input 	int_nxt_addr_reg_dly_3;
input 	int_nxt_addr_reg_dly_2;
input 	clk_clk;
input 	tick_out_external_connection_export;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_mux_out~combout ;


dffeas \readdata[0] (
	.clk(clk_clk),
	.d(\read_mux_out~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

cyclonev_lcell_comb read_mux_out(
	.dataa(!tick_out_external_connection_export),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam read_mux_out.extended_lut = "off";
defparam read_mux_out.lut_mask = 64'h4040404040404040;
defparam read_mux_out.shared_arith = "off";

endmodule

module spw_babasu_spw_babasu_RX_EMPTY_2 (
	altera_reset_synchronizer_int_chain_out,
	readdata_0,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	clk_clk,
	tx_full_external_connection_export)/* synthesis synthesis_greybox=0 */;
input 	altera_reset_synchronizer_int_chain_out;
output 	readdata_0;
input 	int_nxt_addr_reg_dly_3;
input 	int_nxt_addr_reg_dly_2;
input 	clk_clk;
input 	tx_full_external_connection_export;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_mux_out~combout ;


dffeas \readdata[0] (
	.clk(clk_clk),
	.d(\read_mux_out~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

cyclonev_lcell_comb read_mux_out(
	.dataa(!tx_full_external_connection_export),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam read_mux_out.extended_lut = "off";
defparam read_mux_out.lut_mask = 64'h4040404040404040;
defparam read_mux_out.shared_arith = "off";

endmodule

module spw_babasu_spw_babasu_TIME_IN (
	data_out_0,
	data_out_1,
	data_out_2,
	data_out_3,
	data_out_4,
	data_out_5,
	data_out_6,
	data_out_7,
	wait_latency_counter_1,
	wait_latency_counter_0,
	reset_n,
	writedata,
	m0_write,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	readdata_4,
	readdata_5,
	readdata_6,
	readdata_7,
	clk)/* synthesis synthesis_greybox=0 */;
output 	data_out_0;
output 	data_out_1;
output 	data_out_2;
output 	data_out_3;
output 	data_out_4;
output 	data_out_5;
output 	data_out_6;
output 	data_out_7;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	reset_n;
input 	[31:0] writedata;
input 	m0_write;
input 	int_nxt_addr_reg_dly_3;
input 	int_nxt_addr_reg_dly_2;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
output 	readdata_4;
output 	readdata_5;
output 	readdata_6;
output 	readdata_7;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always0~0_combout ;


dffeas \data_out[0] (
	.clk(clk),
	.d(writedata[0]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_0),
	.prn(vcc));
defparam \data_out[0] .is_wysiwyg = "true";
defparam \data_out[0] .power_up = "low";

dffeas \data_out[1] (
	.clk(clk),
	.d(writedata[1]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_1),
	.prn(vcc));
defparam \data_out[1] .is_wysiwyg = "true";
defparam \data_out[1] .power_up = "low";

dffeas \data_out[2] (
	.clk(clk),
	.d(writedata[2]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_2),
	.prn(vcc));
defparam \data_out[2] .is_wysiwyg = "true";
defparam \data_out[2] .power_up = "low";

dffeas \data_out[3] (
	.clk(clk),
	.d(writedata[3]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_3),
	.prn(vcc));
defparam \data_out[3] .is_wysiwyg = "true";
defparam \data_out[3] .power_up = "low";

dffeas \data_out[4] (
	.clk(clk),
	.d(writedata[4]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_4),
	.prn(vcc));
defparam \data_out[4] .is_wysiwyg = "true";
defparam \data_out[4] .power_up = "low";

dffeas \data_out[5] (
	.clk(clk),
	.d(writedata[5]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_5),
	.prn(vcc));
defparam \data_out[5] .is_wysiwyg = "true";
defparam \data_out[5] .power_up = "low";

dffeas \data_out[6] (
	.clk(clk),
	.d(writedata[6]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_6),
	.prn(vcc));
defparam \data_out[6] .is_wysiwyg = "true";
defparam \data_out[6] .power_up = "low";

dffeas \data_out[7] (
	.clk(clk),
	.d(writedata[7]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_7),
	.prn(vcc));
defparam \data_out[7] .is_wysiwyg = "true";
defparam \data_out[7] .power_up = "low";

cyclonev_lcell_comb \readdata[0] (
	.dataa(!data_out_0),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[0] .extended_lut = "off";
defparam \readdata[0] .lut_mask = 64'h4040404040404040;
defparam \readdata[0] .shared_arith = "off";

cyclonev_lcell_comb \readdata[1] (
	.dataa(!data_out_1),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[1] .extended_lut = "off";
defparam \readdata[1] .lut_mask = 64'h4040404040404040;
defparam \readdata[1] .shared_arith = "off";

cyclonev_lcell_comb \readdata[2] (
	.dataa(!data_out_2),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[2] .extended_lut = "off";
defparam \readdata[2] .lut_mask = 64'h4040404040404040;
defparam \readdata[2] .shared_arith = "off";

cyclonev_lcell_comb \readdata[3] (
	.dataa(!data_out_3),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[3] .extended_lut = "off";
defparam \readdata[3] .lut_mask = 64'h4040404040404040;
defparam \readdata[3] .shared_arith = "off";

cyclonev_lcell_comb \readdata[4] (
	.dataa(!data_out_4),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[4] .extended_lut = "off";
defparam \readdata[4] .lut_mask = 64'h4040404040404040;
defparam \readdata[4] .shared_arith = "off";

cyclonev_lcell_comb \readdata[5] (
	.dataa(!data_out_5),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[5] .extended_lut = "off";
defparam \readdata[5] .lut_mask = 64'h4040404040404040;
defparam \readdata[5] .shared_arith = "off";

cyclonev_lcell_comb \readdata[6] (
	.dataa(!data_out_6),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_6),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[6] .extended_lut = "off";
defparam \readdata[6] .lut_mask = 64'h4040404040404040;
defparam \readdata[6] .shared_arith = "off";

cyclonev_lcell_comb \readdata[7] (
	.dataa(!data_out_7),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_7),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[7] .extended_lut = "off";
defparam \readdata[7] .lut_mask = 64'h4040404040404040;
defparam \readdata[7] .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!m0_write),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(!int_nxt_addr_reg_dly_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'h0800000008000000;
defparam \always0~0 .shared_arith = "off";

endmodule

module spw_babasu_spw_babasu_TIME_OUT (
	altera_reset_synchronizer_int_chain_out,
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	readdata_4,
	readdata_5,
	readdata_6,
	readdata_7,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	clk_clk,
	time_out_external_connection_export_0,
	time_out_external_connection_export_1,
	time_out_external_connection_export_2,
	time_out_external_connection_export_3,
	time_out_external_connection_export_4,
	time_out_external_connection_export_5,
	time_out_external_connection_export_6,
	time_out_external_connection_export_7)/* synthesis synthesis_greybox=0 */;
input 	altera_reset_synchronizer_int_chain_out;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
output 	readdata_4;
output 	readdata_5;
output 	readdata_6;
output 	readdata_7;
input 	int_nxt_addr_reg_dly_3;
input 	int_nxt_addr_reg_dly_2;
input 	clk_clk;
input 	time_out_external_connection_export_0;
input 	time_out_external_connection_export_1;
input 	time_out_external_connection_export_2;
input 	time_out_external_connection_export_3;
input 	time_out_external_connection_export_4;
input 	time_out_external_connection_export_5;
input 	time_out_external_connection_export_6;
input 	time_out_external_connection_export_7;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_mux_out[0]~combout ;
wire \read_mux_out[1]~combout ;
wire \read_mux_out[2]~combout ;
wire \read_mux_out[3]~combout ;
wire \read_mux_out[4]~combout ;
wire \read_mux_out[5]~combout ;
wire \read_mux_out[6]~combout ;
wire \read_mux_out[7]~combout ;


dffeas \readdata[0] (
	.clk(clk_clk),
	.d(\read_mux_out[0]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

dffeas \readdata[1] (
	.clk(clk_clk),
	.d(\read_mux_out[1]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_1),
	.prn(vcc));
defparam \readdata[1] .is_wysiwyg = "true";
defparam \readdata[1] .power_up = "low";

dffeas \readdata[2] (
	.clk(clk_clk),
	.d(\read_mux_out[2]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_2),
	.prn(vcc));
defparam \readdata[2] .is_wysiwyg = "true";
defparam \readdata[2] .power_up = "low";

dffeas \readdata[3] (
	.clk(clk_clk),
	.d(\read_mux_out[3]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_3),
	.prn(vcc));
defparam \readdata[3] .is_wysiwyg = "true";
defparam \readdata[3] .power_up = "low";

dffeas \readdata[4] (
	.clk(clk_clk),
	.d(\read_mux_out[4]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_4),
	.prn(vcc));
defparam \readdata[4] .is_wysiwyg = "true";
defparam \readdata[4] .power_up = "low";

dffeas \readdata[5] (
	.clk(clk_clk),
	.d(\read_mux_out[5]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_5),
	.prn(vcc));
defparam \readdata[5] .is_wysiwyg = "true";
defparam \readdata[5] .power_up = "low";

dffeas \readdata[6] (
	.clk(clk_clk),
	.d(\read_mux_out[6]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_6),
	.prn(vcc));
defparam \readdata[6] .is_wysiwyg = "true";
defparam \readdata[6] .power_up = "low";

dffeas \readdata[7] (
	.clk(clk_clk),
	.d(\read_mux_out[7]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_7),
	.prn(vcc));
defparam \readdata[7] .is_wysiwyg = "true";
defparam \readdata[7] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[0] (
	.dataa(!time_out_external_connection_export_0),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[0] .extended_lut = "off";
defparam \read_mux_out[0] .lut_mask = 64'h4040404040404040;
defparam \read_mux_out[0] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[1] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!time_out_external_connection_export_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[1] .extended_lut = "off";
defparam \read_mux_out[1] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[1] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[2] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!time_out_external_connection_export_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[2] .extended_lut = "off";
defparam \read_mux_out[2] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[2] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[3] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!time_out_external_connection_export_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[3] .extended_lut = "off";
defparam \read_mux_out[3] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[3] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[4] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!time_out_external_connection_export_4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[4]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[4] .extended_lut = "off";
defparam \read_mux_out[4] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[4] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[5] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!time_out_external_connection_export_5),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[5]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[5] .extended_lut = "off";
defparam \read_mux_out[5] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[5] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[6] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!time_out_external_connection_export_6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[6]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[6] .extended_lut = "off";
defparam \read_mux_out[6] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[6] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[7] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!time_out_external_connection_export_7),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[7]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[7] .extended_lut = "off";
defparam \read_mux_out[7] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[7] .shared_arith = "off";

endmodule

module spw_babasu_spw_babasu_TX_CLK_DIV (
	data_out_0,
	data_out_1,
	data_out_2,
	data_out_3,
	data_out_4,
	data_out_5,
	data_out_6,
	wait_latency_counter_1,
	wait_latency_counter_0,
	reset_n,
	in_data_reg_0,
	m0_write,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	in_data_reg_1,
	writedata,
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	readdata_4,
	readdata_5,
	readdata_6,
	clk)/* synthesis synthesis_greybox=0 */;
output 	data_out_0;
output 	data_out_1;
output 	data_out_2;
output 	data_out_3;
output 	data_out_4;
output 	data_out_5;
output 	data_out_6;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	reset_n;
input 	in_data_reg_0;
input 	m0_write;
input 	int_nxt_addr_reg_dly_3;
input 	int_nxt_addr_reg_dly_2;
input 	in_data_reg_1;
input 	[31:0] writedata;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
output 	readdata_4;
output 	readdata_5;
output 	readdata_6;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \data_out[0]~0_combout ;
wire \always0~0_combout ;
wire \data_out[1]~1_combout ;


dffeas \data_out[0] (
	.clk(clk),
	.d(\data_out[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_0),
	.prn(vcc));
defparam \data_out[0] .is_wysiwyg = "true";
defparam \data_out[0] .power_up = "low";

dffeas \data_out[1] (
	.clk(clk),
	.d(\data_out[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_1),
	.prn(vcc));
defparam \data_out[1] .is_wysiwyg = "true";
defparam \data_out[1] .power_up = "low";

dffeas \data_out[2] (
	.clk(clk),
	.d(writedata[2]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_2),
	.prn(vcc));
defparam \data_out[2] .is_wysiwyg = "true";
defparam \data_out[2] .power_up = "low";

dffeas \data_out[3] (
	.clk(clk),
	.d(writedata[3]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_3),
	.prn(vcc));
defparam \data_out[3] .is_wysiwyg = "true";
defparam \data_out[3] .power_up = "low";

dffeas \data_out[4] (
	.clk(clk),
	.d(writedata[4]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_4),
	.prn(vcc));
defparam \data_out[4] .is_wysiwyg = "true";
defparam \data_out[4] .power_up = "low";

dffeas \data_out[5] (
	.clk(clk),
	.d(writedata[5]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_5),
	.prn(vcc));
defparam \data_out[5] .is_wysiwyg = "true";
defparam \data_out[5] .power_up = "low";

dffeas \data_out[6] (
	.clk(clk),
	.d(writedata[6]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_6),
	.prn(vcc));
defparam \data_out[6] .is_wysiwyg = "true";
defparam \data_out[6] .power_up = "low";

cyclonev_lcell_comb \readdata[0] (
	.dataa(!data_out_0),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[0] .extended_lut = "off";
defparam \readdata[0] .lut_mask = 64'h8080808080808080;
defparam \readdata[0] .shared_arith = "off";

cyclonev_lcell_comb \readdata[1] (
	.dataa(!data_out_1),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[1] .extended_lut = "off";
defparam \readdata[1] .lut_mask = 64'h8080808080808080;
defparam \readdata[1] .shared_arith = "off";

cyclonev_lcell_comb \readdata[2] (
	.dataa(!data_out_2),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[2] .extended_lut = "off";
defparam \readdata[2] .lut_mask = 64'h4040404040404040;
defparam \readdata[2] .shared_arith = "off";

cyclonev_lcell_comb \readdata[3] (
	.dataa(!data_out_3),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[3] .extended_lut = "off";
defparam \readdata[3] .lut_mask = 64'h4040404040404040;
defparam \readdata[3] .shared_arith = "off";

cyclonev_lcell_comb \readdata[4] (
	.dataa(!data_out_4),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[4] .extended_lut = "off";
defparam \readdata[4] .lut_mask = 64'h4040404040404040;
defparam \readdata[4] .shared_arith = "off";

cyclonev_lcell_comb \readdata[5] (
	.dataa(!data_out_5),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[5] .extended_lut = "off";
defparam \readdata[5] .lut_mask = 64'h4040404040404040;
defparam \readdata[5] .shared_arith = "off";

cyclonev_lcell_comb \readdata[6] (
	.dataa(!data_out_6),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_6),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[6] .extended_lut = "off";
defparam \readdata[6] .lut_mask = 64'h4040404040404040;
defparam \readdata[6] .shared_arith = "off";

cyclonev_lcell_comb \data_out[0]~0 (
	.dataa(!in_data_reg_0),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out[0]~0 .extended_lut = "off";
defparam \data_out[0]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \data_out[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!m0_write),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(!int_nxt_addr_reg_dly_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'h0800000008000000;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \data_out[1]~1 (
	.dataa(!in_data_reg_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out[1]~1 .extended_lut = "off";
defparam \data_out[1]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \data_out[1]~1 .shared_arith = "off";

endmodule
