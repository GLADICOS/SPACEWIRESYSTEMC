// jaxa.v

// Generated using ACDS version 17.1 593

`timescale 1 ps / 1 ps
module jaxa (
		output wire        autostart_external_connection_export,                   //                   autostart_external_connection.export
		input  wire        clk_clk,                                                //                                             clk.clk
		output wire [1:0]  controlflagsin_external_connection_export,              //              controlflagsin_external_connection.export
		input  wire [1:0]  controlflagsout_external_connection_export,             //             controlflagsout_external_connection.export
		input  wire [5:0]  creditcount_external_connection_export,                 //                 creditcount_external_connection.export
		input  wire [7:0]  errorstatus_external_connection_export,                 //                 errorstatus_external_connection.export
		output wire        linkdisable_external_connection_export,                 //                 linkdisable_external_connection.export
		output wire        linkstart_external_connection_export,                   //                   linkstart_external_connection.export
		input  wire [15:0] linkstatus_external_connection_export,                  //                  linkstatus_external_connection.export
		output wire [12:0] memory_mem_a,                                           //                                          memory.mem_a
		output wire [2:0]  memory_mem_ba,                                          //                                                .mem_ba
		output wire        memory_mem_ck,                                          //                                                .mem_ck
		output wire        memory_mem_ck_n,                                        //                                                .mem_ck_n
		output wire        memory_mem_cke,                                         //                                                .mem_cke
		output wire        memory_mem_cs_n,                                        //                                                .mem_cs_n
		output wire        memory_mem_ras_n,                                       //                                                .mem_ras_n
		output wire        memory_mem_cas_n,                                       //                                                .mem_cas_n
		output wire        memory_mem_we_n,                                        //                                                .mem_we_n
		output wire        memory_mem_reset_n,                                     //                                                .mem_reset_n
		inout  wire [7:0]  memory_mem_dq,                                          //                                                .mem_dq
		inout  wire        memory_mem_dqs,                                         //                                                .mem_dqs
		inout  wire        memory_mem_dqs_n,                                       //                                                .mem_dqs_n
		output wire        memory_mem_odt,                                         //                                                .mem_odt
		output wire        memory_mem_dm,                                          //                                                .mem_dm
		input  wire        memory_oct_rzqin,                                       //                                                .oct_rzqin
		input  wire [5:0]  outstandingcount_external_connection_export,            //            outstandingcount_external_connection.export
		output wire        pll_0_outclk0_clk,                                      //                                   pll_0_outclk0.clk
		input  wire        receiveactivity_external_connection_export,             //             receiveactivity_external_connection.export
		output wire        receiveclock_external_connection_export,                //                receiveclock_external_connection.export
		input  wire        receivefifodatacount_external_connection_export,        //        receivefifodatacount_external_connection.export
		input  wire [8:0]  receivefifodataout_external_connection_export,          //          receivefifodataout_external_connection.export
		input  wire        receivefifoempty_external_connection_export,            //            receivefifoempty_external_connection.export
		input  wire        receivefifofull_external_connection_export,             //             receivefifofull_external_connection.export
		output wire        receivefiforeadenable_external_connection_export,       //       receivefiforeadenable_external_connection.export
		output wire        spacewiredatain_external_connection_export,             //             spacewiredatain_external_connection.export
		input  wire        spacewiredataout_external_connection_export,            //            spacewiredataout_external_connection.export
		output wire        spacewirestrobein_external_connection_export,           //           spacewirestrobein_external_connection.export
		input  wire        spacewirestrobeout_external_connection_export,          //          spacewirestrobeout_external_connection.export
		input  wire [31:0] statisticalinformation_0_external_connection_export,    //    statisticalinformation_0_external_connection.export
		output wire [7:0]  statisticalinformation_1_external_connection_export,    //    statisticalinformation_1_external_connection.export
		output wire        statisticalinformationclear_external_connection_export, // statisticalinformationclear_external_connection.export
		output wire        tickin_external_connection_export,                      //                      tickin_external_connection.export
		input  wire        tickout_external_connection_export,                     //                     tickout_external_connection.export
		output wire [5:0]  timein_external_connection_export,                      //                      timein_external_connection.export
		input  wire [5:0]  timeout_external_connection_export,                     //                     timeout_external_connection.export
		input  wire        transmitactivity_external_connection_export,            //            transmitactivity_external_connection.export
		output wire        transmitclock_external_connection_export,               //               transmitclock_external_connection.export
		output wire [5:0]  transmitclockdividevalue_external_connection_export,    //    transmitclockdividevalue_external_connection.export
		input  wire [5:0]  transmitfifodatacount_external_connection_export,       //       transmitfifodatacount_external_connection.export
		output wire [8:0]  transmitfifodatain_external_connection_export,          //          transmitfifodatain_external_connection.export
		input  wire        transmitfifofull_external_connection_export,            //            transmitfifofull_external_connection.export
		output wire        transmitfifowriteenable_external_connection_export      //     transmitfifowriteenable_external_connection.export
	);

	wire         hps_0_h2f_reset_reset;                                       // hps_0:h2f_rst_n -> [pll_0:rst, rst_controller:reset_in0, rst_controller_001:reset_in0]
	wire   [1:0] hps_0_h2f_axi_master_awburst;                                // hps_0:h2f_AWBURST -> mm_interconnect_0:hps_0_h2f_axi_master_awburst
	wire   [3:0] hps_0_h2f_axi_master_arlen;                                  // hps_0:h2f_ARLEN -> mm_interconnect_0:hps_0_h2f_axi_master_arlen
	wire   [3:0] hps_0_h2f_axi_master_wstrb;                                  // hps_0:h2f_WSTRB -> mm_interconnect_0:hps_0_h2f_axi_master_wstrb
	wire         hps_0_h2f_axi_master_wready;                                 // mm_interconnect_0:hps_0_h2f_axi_master_wready -> hps_0:h2f_WREADY
	wire  [11:0] hps_0_h2f_axi_master_rid;                                    // mm_interconnect_0:hps_0_h2f_axi_master_rid -> hps_0:h2f_RID
	wire         hps_0_h2f_axi_master_rready;                                 // hps_0:h2f_RREADY -> mm_interconnect_0:hps_0_h2f_axi_master_rready
	wire   [3:0] hps_0_h2f_axi_master_awlen;                                  // hps_0:h2f_AWLEN -> mm_interconnect_0:hps_0_h2f_axi_master_awlen
	wire  [11:0] hps_0_h2f_axi_master_wid;                                    // hps_0:h2f_WID -> mm_interconnect_0:hps_0_h2f_axi_master_wid
	wire   [3:0] hps_0_h2f_axi_master_arcache;                                // hps_0:h2f_ARCACHE -> mm_interconnect_0:hps_0_h2f_axi_master_arcache
	wire         hps_0_h2f_axi_master_wvalid;                                 // hps_0:h2f_WVALID -> mm_interconnect_0:hps_0_h2f_axi_master_wvalid
	wire  [29:0] hps_0_h2f_axi_master_araddr;                                 // hps_0:h2f_ARADDR -> mm_interconnect_0:hps_0_h2f_axi_master_araddr
	wire   [2:0] hps_0_h2f_axi_master_arprot;                                 // hps_0:h2f_ARPROT -> mm_interconnect_0:hps_0_h2f_axi_master_arprot
	wire   [2:0] hps_0_h2f_axi_master_awprot;                                 // hps_0:h2f_AWPROT -> mm_interconnect_0:hps_0_h2f_axi_master_awprot
	wire  [31:0] hps_0_h2f_axi_master_wdata;                                  // hps_0:h2f_WDATA -> mm_interconnect_0:hps_0_h2f_axi_master_wdata
	wire         hps_0_h2f_axi_master_arvalid;                                // hps_0:h2f_ARVALID -> mm_interconnect_0:hps_0_h2f_axi_master_arvalid
	wire   [3:0] hps_0_h2f_axi_master_awcache;                                // hps_0:h2f_AWCACHE -> mm_interconnect_0:hps_0_h2f_axi_master_awcache
	wire  [11:0] hps_0_h2f_axi_master_arid;                                   // hps_0:h2f_ARID -> mm_interconnect_0:hps_0_h2f_axi_master_arid
	wire   [1:0] hps_0_h2f_axi_master_arlock;                                 // hps_0:h2f_ARLOCK -> mm_interconnect_0:hps_0_h2f_axi_master_arlock
	wire   [1:0] hps_0_h2f_axi_master_awlock;                                 // hps_0:h2f_AWLOCK -> mm_interconnect_0:hps_0_h2f_axi_master_awlock
	wire  [29:0] hps_0_h2f_axi_master_awaddr;                                 // hps_0:h2f_AWADDR -> mm_interconnect_0:hps_0_h2f_axi_master_awaddr
	wire   [1:0] hps_0_h2f_axi_master_bresp;                                  // mm_interconnect_0:hps_0_h2f_axi_master_bresp -> hps_0:h2f_BRESP
	wire         hps_0_h2f_axi_master_arready;                                // mm_interconnect_0:hps_0_h2f_axi_master_arready -> hps_0:h2f_ARREADY
	wire  [31:0] hps_0_h2f_axi_master_rdata;                                  // mm_interconnect_0:hps_0_h2f_axi_master_rdata -> hps_0:h2f_RDATA
	wire         hps_0_h2f_axi_master_awready;                                // mm_interconnect_0:hps_0_h2f_axi_master_awready -> hps_0:h2f_AWREADY
	wire   [1:0] hps_0_h2f_axi_master_arburst;                                // hps_0:h2f_ARBURST -> mm_interconnect_0:hps_0_h2f_axi_master_arburst
	wire   [2:0] hps_0_h2f_axi_master_arsize;                                 // hps_0:h2f_ARSIZE -> mm_interconnect_0:hps_0_h2f_axi_master_arsize
	wire         hps_0_h2f_axi_master_bready;                                 // hps_0:h2f_BREADY -> mm_interconnect_0:hps_0_h2f_axi_master_bready
	wire         hps_0_h2f_axi_master_rlast;                                  // mm_interconnect_0:hps_0_h2f_axi_master_rlast -> hps_0:h2f_RLAST
	wire         hps_0_h2f_axi_master_wlast;                                  // hps_0:h2f_WLAST -> mm_interconnect_0:hps_0_h2f_axi_master_wlast
	wire   [1:0] hps_0_h2f_axi_master_rresp;                                  // mm_interconnect_0:hps_0_h2f_axi_master_rresp -> hps_0:h2f_RRESP
	wire  [11:0] hps_0_h2f_axi_master_awid;                                   // hps_0:h2f_AWID -> mm_interconnect_0:hps_0_h2f_axi_master_awid
	wire  [11:0] hps_0_h2f_axi_master_bid;                                    // mm_interconnect_0:hps_0_h2f_axi_master_bid -> hps_0:h2f_BID
	wire         hps_0_h2f_axi_master_bvalid;                                 // mm_interconnect_0:hps_0_h2f_axi_master_bvalid -> hps_0:h2f_BVALID
	wire   [2:0] hps_0_h2f_axi_master_awsize;                                 // hps_0:h2f_AWSIZE -> mm_interconnect_0:hps_0_h2f_axi_master_awsize
	wire         hps_0_h2f_axi_master_awvalid;                                // hps_0:h2f_AWVALID -> mm_interconnect_0:hps_0_h2f_axi_master_awvalid
	wire         hps_0_h2f_axi_master_rvalid;                                 // mm_interconnect_0:hps_0_h2f_axi_master_rvalid -> hps_0:h2f_RVALID
	wire         mm_interconnect_0_autostart_s1_chipselect;                   // mm_interconnect_0:autoStart_s1_chipselect -> autoStart:chipselect
	wire  [31:0] mm_interconnect_0_autostart_s1_readdata;                     // autoStart:readdata -> mm_interconnect_0:autoStart_s1_readdata
	wire   [1:0] mm_interconnect_0_autostart_s1_address;                      // mm_interconnect_0:autoStart_s1_address -> autoStart:address
	wire         mm_interconnect_0_autostart_s1_write;                        // mm_interconnect_0:autoStart_s1_write -> autoStart:write_n
	wire  [31:0] mm_interconnect_0_autostart_s1_writedata;                    // mm_interconnect_0:autoStart_s1_writedata -> autoStart:writedata
	wire         mm_interconnect_0_linkdisable_s1_chipselect;                 // mm_interconnect_0:linkDisable_s1_chipselect -> linkDisable:chipselect
	wire  [31:0] mm_interconnect_0_linkdisable_s1_readdata;                   // linkDisable:readdata -> mm_interconnect_0:linkDisable_s1_readdata
	wire   [1:0] mm_interconnect_0_linkdisable_s1_address;                    // mm_interconnect_0:linkDisable_s1_address -> linkDisable:address
	wire         mm_interconnect_0_linkdisable_s1_write;                      // mm_interconnect_0:linkDisable_s1_write -> linkDisable:write_n
	wire  [31:0] mm_interconnect_0_linkdisable_s1_writedata;                  // mm_interconnect_0:linkDisable_s1_writedata -> linkDisable:writedata
	wire         mm_interconnect_0_linkstart_s1_chipselect;                   // mm_interconnect_0:linkStart_s1_chipselect -> linkStart:chipselect
	wire  [31:0] mm_interconnect_0_linkstart_s1_readdata;                     // linkStart:readdata -> mm_interconnect_0:linkStart_s1_readdata
	wire   [1:0] mm_interconnect_0_linkstart_s1_address;                      // mm_interconnect_0:linkStart_s1_address -> linkStart:address
	wire         mm_interconnect_0_linkstart_s1_write;                        // mm_interconnect_0:linkStart_s1_write -> linkStart:write_n
	wire  [31:0] mm_interconnect_0_linkstart_s1_writedata;                    // mm_interconnect_0:linkStart_s1_writedata -> linkStart:writedata
	wire  [31:0] mm_interconnect_0_receivefifodatacount_s1_readdata;          // receiveFIFODataCount:readdata -> mm_interconnect_0:receiveFIFODataCount_s1_readdata
	wire   [1:0] mm_interconnect_0_receivefifodatacount_s1_address;           // mm_interconnect_0:receiveFIFODataCount_s1_address -> receiveFIFODataCount:address
	wire  [31:0] mm_interconnect_0_receivefifodataout_s1_readdata;            // receiveFIFODataOut:readdata -> mm_interconnect_0:receiveFIFODataOut_s1_readdata
	wire   [1:0] mm_interconnect_0_receivefifodataout_s1_address;             // mm_interconnect_0:receiveFIFODataOut_s1_address -> receiveFIFODataOut:address
	wire  [31:0] mm_interconnect_0_receivefifoempty_s1_readdata;              // receiveFIFOEmpty:readdata -> mm_interconnect_0:receiveFIFOEmpty_s1_readdata
	wire   [1:0] mm_interconnect_0_receivefifoempty_s1_address;               // mm_interconnect_0:receiveFIFOEmpty_s1_address -> receiveFIFOEmpty:address
	wire  [31:0] mm_interconnect_0_receivefifofull_s1_readdata;               // receiveFIFOFull:readdata -> mm_interconnect_0:receiveFIFOFull_s1_readdata
	wire   [1:0] mm_interconnect_0_receivefifofull_s1_address;                // mm_interconnect_0:receiveFIFOFull_s1_address -> receiveFIFOFull:address
	wire         mm_interconnect_0_receivefiforeadenable_s1_chipselect;       // mm_interconnect_0:receiveFIFOReadEnable_s1_chipselect -> receiveFIFOReadEnable:chipselect
	wire  [31:0] mm_interconnect_0_receivefiforeadenable_s1_readdata;         // receiveFIFOReadEnable:readdata -> mm_interconnect_0:receiveFIFOReadEnable_s1_readdata
	wire   [1:0] mm_interconnect_0_receivefiforeadenable_s1_address;          // mm_interconnect_0:receiveFIFOReadEnable_s1_address -> receiveFIFOReadEnable:address
	wire         mm_interconnect_0_receivefiforeadenable_s1_write;            // mm_interconnect_0:receiveFIFOReadEnable_s1_write -> receiveFIFOReadEnable:write_n
	wire  [31:0] mm_interconnect_0_receivefiforeadenable_s1_writedata;        // mm_interconnect_0:receiveFIFOReadEnable_s1_writedata -> receiveFIFOReadEnable:writedata
	wire  [31:0] mm_interconnect_0_transmitfifofull_s1_readdata;              // transmitFIFOFull:readdata -> mm_interconnect_0:transmitFIFOFull_s1_readdata
	wire   [1:0] mm_interconnect_0_transmitfifofull_s1_address;               // mm_interconnect_0:transmitFIFOFull_s1_address -> transmitFIFOFull:address
	wire         mm_interconnect_0_transmitfifowriteenable_s1_chipselect;     // mm_interconnect_0:transmitFIFOWriteEnable_s1_chipselect -> transmitFIFOWriteEnable:chipselect
	wire  [31:0] mm_interconnect_0_transmitfifowriteenable_s1_readdata;       // transmitFIFOWriteEnable:readdata -> mm_interconnect_0:transmitFIFOWriteEnable_s1_readdata
	wire   [1:0] mm_interconnect_0_transmitfifowriteenable_s1_address;        // mm_interconnect_0:transmitFIFOWriteEnable_s1_address -> transmitFIFOWriteEnable:address
	wire         mm_interconnect_0_transmitfifowriteenable_s1_write;          // mm_interconnect_0:transmitFIFOWriteEnable_s1_write -> transmitFIFOWriteEnable:write_n
	wire  [31:0] mm_interconnect_0_transmitfifowriteenable_s1_writedata;      // mm_interconnect_0:transmitFIFOWriteEnable_s1_writedata -> transmitFIFOWriteEnable:writedata
	wire         mm_interconnect_0_transmitfifodatain_s1_chipselect;          // mm_interconnect_0:transmitFIFODataIn_s1_chipselect -> transmitFIFODataIn:chipselect
	wire  [31:0] mm_interconnect_0_transmitfifodatain_s1_readdata;            // transmitFIFODataIn:readdata -> mm_interconnect_0:transmitFIFODataIn_s1_readdata
	wire   [1:0] mm_interconnect_0_transmitfifodatain_s1_address;             // mm_interconnect_0:transmitFIFODataIn_s1_address -> transmitFIFODataIn:address
	wire         mm_interconnect_0_transmitfifodatain_s1_write;               // mm_interconnect_0:transmitFIFODataIn_s1_write -> transmitFIFODataIn:write_n
	wire  [31:0] mm_interconnect_0_transmitfifodatain_s1_writedata;           // mm_interconnect_0:transmitFIFODataIn_s1_writedata -> transmitFIFODataIn:writedata
	wire  [31:0] mm_interconnect_0_transmitfifodatacount_s1_readdata;         // transmitFIFODataCount:readdata -> mm_interconnect_0:transmitFIFODataCount_s1_readdata
	wire   [1:0] mm_interconnect_0_transmitfifodatacount_s1_address;          // mm_interconnect_0:transmitFIFODataCount_s1_address -> transmitFIFODataCount:address
	wire         mm_interconnect_0_tickin_s1_chipselect;                      // mm_interconnect_0:tickIn_s1_chipselect -> tickIn:chipselect
	wire  [31:0] mm_interconnect_0_tickin_s1_readdata;                        // tickIn:readdata -> mm_interconnect_0:tickIn_s1_readdata
	wire   [1:0] mm_interconnect_0_tickin_s1_address;                         // mm_interconnect_0:tickIn_s1_address -> tickIn:address
	wire         mm_interconnect_0_tickin_s1_write;                           // mm_interconnect_0:tickIn_s1_write -> tickIn:write_n
	wire  [31:0] mm_interconnect_0_tickin_s1_writedata;                       // mm_interconnect_0:tickIn_s1_writedata -> tickIn:writedata
	wire         mm_interconnect_0_timein_s1_chipselect;                      // mm_interconnect_0:timeIn_s1_chipselect -> timeIn:chipselect
	wire  [31:0] mm_interconnect_0_timein_s1_readdata;                        // timeIn:readdata -> mm_interconnect_0:timeIn_s1_readdata
	wire   [1:0] mm_interconnect_0_timein_s1_address;                         // mm_interconnect_0:timeIn_s1_address -> timeIn:address
	wire         mm_interconnect_0_timein_s1_write;                           // mm_interconnect_0:timeIn_s1_write -> timeIn:write_n
	wire  [31:0] mm_interconnect_0_timein_s1_writedata;                       // mm_interconnect_0:timeIn_s1_writedata -> timeIn:writedata
	wire  [31:0] mm_interconnect_0_tickout_s1_readdata;                       // tickOut:readdata -> mm_interconnect_0:tickOut_s1_readdata
	wire   [1:0] mm_interconnect_0_tickout_s1_address;                        // mm_interconnect_0:tickOut_s1_address -> tickOut:address
	wire  [31:0] mm_interconnect_0_timeout_s1_readdata;                       // timeOut:readdata -> mm_interconnect_0:timeOut_s1_readdata
	wire   [1:0] mm_interconnect_0_timeout_s1_address;                        // mm_interconnect_0:timeOut_s1_address -> timeOut:address
	wire  [31:0] mm_interconnect_0_statisticalinformation_0_s1_readdata;      // statisticalInformation_0:readdata -> mm_interconnect_0:statisticalInformation_0_s1_readdata
	wire   [1:0] mm_interconnect_0_statisticalinformation_0_s1_address;       // mm_interconnect_0:statisticalInformation_0_s1_address -> statisticalInformation_0:address
	wire         mm_interconnect_0_statisticalinformation_1_s1_chipselect;    // mm_interconnect_0:statisticalInformation_1_s1_chipselect -> statisticalInformation_1:chipselect
	wire  [31:0] mm_interconnect_0_statisticalinformation_1_s1_readdata;      // statisticalInformation_1:readdata -> mm_interconnect_0:statisticalInformation_1_s1_readdata
	wire   [1:0] mm_interconnect_0_statisticalinformation_1_s1_address;       // mm_interconnect_0:statisticalInformation_1_s1_address -> statisticalInformation_1:address
	wire         mm_interconnect_0_statisticalinformation_1_s1_write;         // mm_interconnect_0:statisticalInformation_1_s1_write -> statisticalInformation_1:write_n
	wire  [31:0] mm_interconnect_0_statisticalinformation_1_s1_writedata;     // mm_interconnect_0:statisticalInformation_1_s1_writedata -> statisticalInformation_1:writedata
	wire         mm_interconnect_0_statisticalinformationclear_s1_chipselect; // mm_interconnect_0:statisticalInformationClear_s1_chipselect -> statisticalInformationClear:chipselect
	wire  [31:0] mm_interconnect_0_statisticalinformationclear_s1_readdata;   // statisticalInformationClear:readdata -> mm_interconnect_0:statisticalInformationClear_s1_readdata
	wire   [1:0] mm_interconnect_0_statisticalinformationclear_s1_address;    // mm_interconnect_0:statisticalInformationClear_s1_address -> statisticalInformationClear:address
	wire         mm_interconnect_0_statisticalinformationclear_s1_write;      // mm_interconnect_0:statisticalInformationClear_s1_write -> statisticalInformationClear:write_n
	wire  [31:0] mm_interconnect_0_statisticalinformationclear_s1_writedata;  // mm_interconnect_0:statisticalInformationClear_s1_writedata -> statisticalInformationClear:writedata
	wire  [31:0] mm_interconnect_0_linkstatus_s1_readdata;                    // linkStatus:readdata -> mm_interconnect_0:linkStatus_s1_readdata
	wire   [1:0] mm_interconnect_0_linkstatus_s1_address;                     // mm_interconnect_0:linkStatus_s1_address -> linkStatus:address
	wire  [31:0] mm_interconnect_0_errorstatus_s1_readdata;                   // errorStatus:readdata -> mm_interconnect_0:errorStatus_s1_readdata
	wire   [1:0] mm_interconnect_0_errorstatus_s1_address;                    // mm_interconnect_0:errorStatus_s1_address -> errorStatus:address
	wire         mm_interconnect_0_transmitclockdividevalue_s1_chipselect;    // mm_interconnect_0:transmitClockDivideValue_s1_chipselect -> transmitClockDivideValue:chipselect
	wire  [31:0] mm_interconnect_0_transmitclockdividevalue_s1_readdata;      // transmitClockDivideValue:readdata -> mm_interconnect_0:transmitClockDivideValue_s1_readdata
	wire   [1:0] mm_interconnect_0_transmitclockdividevalue_s1_address;       // mm_interconnect_0:transmitClockDivideValue_s1_address -> transmitClockDivideValue:address
	wire         mm_interconnect_0_transmitclockdividevalue_s1_write;         // mm_interconnect_0:transmitClockDivideValue_s1_write -> transmitClockDivideValue:write_n
	wire  [31:0] mm_interconnect_0_transmitclockdividevalue_s1_writedata;     // mm_interconnect_0:transmitClockDivideValue_s1_writedata -> transmitClockDivideValue:writedata
	wire         mm_interconnect_0_transmitclock_s1_chipselect;               // mm_interconnect_0:transmitClock_s1_chipselect -> transmitClock:chipselect
	wire  [31:0] mm_interconnect_0_transmitclock_s1_readdata;                 // transmitClock:readdata -> mm_interconnect_0:transmitClock_s1_readdata
	wire   [1:0] mm_interconnect_0_transmitclock_s1_address;                  // mm_interconnect_0:transmitClock_s1_address -> transmitClock:address
	wire         mm_interconnect_0_transmitclock_s1_write;                    // mm_interconnect_0:transmitClock_s1_write -> transmitClock:write_n
	wire  [31:0] mm_interconnect_0_transmitclock_s1_writedata;                // mm_interconnect_0:transmitClock_s1_writedata -> transmitClock:writedata
	wire  [31:0] mm_interconnect_0_transmitactivity_s1_readdata;              // transmitActivity:readdata -> mm_interconnect_0:transmitActivity_s1_readdata
	wire   [1:0] mm_interconnect_0_transmitactivity_s1_address;               // mm_interconnect_0:transmitActivity_s1_address -> transmitActivity:address
	wire         mm_interconnect_0_spacewirestrobein_s1_chipselect;           // mm_interconnect_0:spaceWireStrobeIn_s1_chipselect -> spaceWireStrobeIn:chipselect
	wire  [31:0] mm_interconnect_0_spacewirestrobein_s1_readdata;             // spaceWireStrobeIn:readdata -> mm_interconnect_0:spaceWireStrobeIn_s1_readdata
	wire   [1:0] mm_interconnect_0_spacewirestrobein_s1_address;              // mm_interconnect_0:spaceWireStrobeIn_s1_address -> spaceWireStrobeIn:address
	wire         mm_interconnect_0_spacewirestrobein_s1_write;                // mm_interconnect_0:spaceWireStrobeIn_s1_write -> spaceWireStrobeIn:write_n
	wire  [31:0] mm_interconnect_0_spacewirestrobein_s1_writedata;            // mm_interconnect_0:spaceWireStrobeIn_s1_writedata -> spaceWireStrobeIn:writedata
	wire  [31:0] mm_interconnect_0_spacewirestrobeout_s1_readdata;            // spaceWireStrobeOut:readdata -> mm_interconnect_0:spaceWireStrobeOut_s1_readdata
	wire   [1:0] mm_interconnect_0_spacewirestrobeout_s1_address;             // mm_interconnect_0:spaceWireStrobeOut_s1_address -> spaceWireStrobeOut:address
	wire  [31:0] mm_interconnect_0_spacewiredataout_s1_readdata;              // spaceWireDataOut:readdata -> mm_interconnect_0:spaceWireDataOut_s1_readdata
	wire   [1:0] mm_interconnect_0_spacewiredataout_s1_address;               // mm_interconnect_0:spaceWireDataOut_s1_address -> spaceWireDataOut:address
	wire         mm_interconnect_0_spacewiredatain_s1_chipselect;             // mm_interconnect_0:spaceWireDataIn_s1_chipselect -> spaceWireDataIn:chipselect
	wire  [31:0] mm_interconnect_0_spacewiredatain_s1_readdata;               // spaceWireDataIn:readdata -> mm_interconnect_0:spaceWireDataIn_s1_readdata
	wire   [1:0] mm_interconnect_0_spacewiredatain_s1_address;                // mm_interconnect_0:spaceWireDataIn_s1_address -> spaceWireDataIn:address
	wire         mm_interconnect_0_spacewiredatain_s1_write;                  // mm_interconnect_0:spaceWireDataIn_s1_write -> spaceWireDataIn:write_n
	wire  [31:0] mm_interconnect_0_spacewiredatain_s1_writedata;              // mm_interconnect_0:spaceWireDataIn_s1_writedata -> spaceWireDataIn:writedata
	wire         mm_interconnect_0_controlflagsin_s1_chipselect;              // mm_interconnect_0:controlFlagsIn_s1_chipselect -> controlFlagsIn:chipselect
	wire  [31:0] mm_interconnect_0_controlflagsin_s1_readdata;                // controlFlagsIn:readdata -> mm_interconnect_0:controlFlagsIn_s1_readdata
	wire   [1:0] mm_interconnect_0_controlflagsin_s1_address;                 // mm_interconnect_0:controlFlagsIn_s1_address -> controlFlagsIn:address
	wire         mm_interconnect_0_controlflagsin_s1_write;                   // mm_interconnect_0:controlFlagsIn_s1_write -> controlFlagsIn:write_n
	wire  [31:0] mm_interconnect_0_controlflagsin_s1_writedata;               // mm_interconnect_0:controlFlagsIn_s1_writedata -> controlFlagsIn:writedata
	wire  [31:0] mm_interconnect_0_controlflagsout_s1_readdata;               // controlFlagsOut:readdata -> mm_interconnect_0:controlFlagsOut_s1_readdata
	wire   [1:0] mm_interconnect_0_controlflagsout_s1_address;                // mm_interconnect_0:controlFlagsOut_s1_address -> controlFlagsOut:address
	wire  [31:0] mm_interconnect_0_creditcount_s1_readdata;                   // creditCount:readdata -> mm_interconnect_0:creditCount_s1_readdata
	wire   [1:0] mm_interconnect_0_creditcount_s1_address;                    // mm_interconnect_0:creditCount_s1_address -> creditCount:address
	wire  [31:0] mm_interconnect_0_outstandingcount_s1_readdata;              // outstandingCount:readdata -> mm_interconnect_0:outstandingCount_s1_readdata
	wire   [1:0] mm_interconnect_0_outstandingcount_s1_address;               // mm_interconnect_0:outstandingCount_s1_address -> outstandingCount:address
	wire  [31:0] mm_interconnect_0_receiveactivity_s1_readdata;               // receiveActivity:readdata -> mm_interconnect_0:receiveActivity_s1_readdata
	wire   [1:0] mm_interconnect_0_receiveactivity_s1_address;                // mm_interconnect_0:receiveActivity_s1_address -> receiveActivity:address
	wire         mm_interconnect_0_receiveclock_s1_chipselect;                // mm_interconnect_0:receiveClock_s1_chipselect -> receiveClock:chipselect
	wire  [31:0] mm_interconnect_0_receiveclock_s1_readdata;                  // receiveClock:readdata -> mm_interconnect_0:receiveClock_s1_readdata
	wire   [1:0] mm_interconnect_0_receiveclock_s1_address;                   // mm_interconnect_0:receiveClock_s1_address -> receiveClock:address
	wire         mm_interconnect_0_receiveclock_s1_write;                     // mm_interconnect_0:receiveClock_s1_write -> receiveClock:write_n
	wire  [31:0] mm_interconnect_0_receiveclock_s1_writedata;                 // mm_interconnect_0:receiveClock_s1_writedata -> receiveClock:writedata
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [autoStart:reset_n, controlFlagsIn:reset_n, controlFlagsOut:reset_n, creditCount:reset_n, errorStatus:reset_n, linkDisable:reset_n, linkStart:reset_n, linkStatus:reset_n, mm_interconnect_0:autoStart_reset_reset_bridge_in_reset_reset, outstandingCount:reset_n, receiveActivity:reset_n, receiveClock:reset_n, receiveFIFODataCount:reset_n, receiveFIFODataOut:reset_n, receiveFIFOEmpty:reset_n, receiveFIFOFull:reset_n, receiveFIFOReadEnable:reset_n, spaceWireDataIn:reset_n, spaceWireDataOut:reset_n, spaceWireStrobeIn:reset_n, spaceWireStrobeOut:reset_n, statisticalInformationClear:reset_n, statisticalInformation_0:reset_n, statisticalInformation_1:reset_n, tickIn:reset_n, tickOut:reset_n, timeIn:reset_n, timeOut:reset_n, transmitActivity:reset_n, transmitClock:reset_n, transmitClockDivideValue:reset_n, transmitFIFODataCount:reset_n, transmitFIFODataIn:reset_n, transmitFIFOFull:reset_n, transmitFIFOWriteEnable:reset_n]
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> mm_interconnect_0:hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset

	jaxa_autoStart autostart (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_autostart_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_autostart_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_autostart_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_autostart_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_autostart_s1_readdata),   //                    .readdata
		.out_port   (autostart_external_connection_export)       // external_connection.export
	);

	jaxa_controlFlagsIn controlflagsin (
		.clk        (clk_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_controlflagsin_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_controlflagsin_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_controlflagsin_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_controlflagsin_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_controlflagsin_s1_readdata),   //                    .readdata
		.out_port   (controlflagsin_external_connection_export)       // external_connection.export
	);

	jaxa_controlFlagsOut controlflagsout (
		.clk      (clk_clk),                                       //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address  (mm_interconnect_0_controlflagsout_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_controlflagsout_s1_readdata), //                    .readdata
		.in_port  (controlflagsout_external_connection_export)     // external_connection.export
	);

	jaxa_creditCount creditcount (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_0_creditcount_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_creditcount_s1_readdata), //                    .readdata
		.in_port  (creditcount_external_connection_export)     // external_connection.export
	);

	jaxa_errorStatus errorstatus (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_0_errorstatus_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_errorstatus_s1_readdata), //                    .readdata
		.in_port  (errorstatus_external_connection_export)     // external_connection.export
	);

	jaxa_hps_0 #(
		.F2S_Width (0),
		.S2F_Width (1)
	) hps_0 (
		.mem_a       (memory_mem_a),                 //         memory.mem_a
		.mem_ba      (memory_mem_ba),                //               .mem_ba
		.mem_ck      (memory_mem_ck),                //               .mem_ck
		.mem_ck_n    (memory_mem_ck_n),              //               .mem_ck_n
		.mem_cke     (memory_mem_cke),               //               .mem_cke
		.mem_cs_n    (memory_mem_cs_n),              //               .mem_cs_n
		.mem_ras_n   (memory_mem_ras_n),             //               .mem_ras_n
		.mem_cas_n   (memory_mem_cas_n),             //               .mem_cas_n
		.mem_we_n    (memory_mem_we_n),              //               .mem_we_n
		.mem_reset_n (memory_mem_reset_n),           //               .mem_reset_n
		.mem_dq      (memory_mem_dq),                //               .mem_dq
		.mem_dqs     (memory_mem_dqs),               //               .mem_dqs
		.mem_dqs_n   (memory_mem_dqs_n),             //               .mem_dqs_n
		.mem_odt     (memory_mem_odt),               //               .mem_odt
		.mem_dm      (memory_mem_dm),                //               .mem_dm
		.oct_rzqin   (memory_oct_rzqin),             //               .oct_rzqin
		.h2f_rst_n   (hps_0_h2f_reset_reset),        //      h2f_reset.reset_n
		.h2f_axi_clk (clk_clk),                      //  h2f_axi_clock.clk
		.h2f_AWID    (hps_0_h2f_axi_master_awid),    // h2f_axi_master.awid
		.h2f_AWADDR  (hps_0_h2f_axi_master_awaddr),  //               .awaddr
		.h2f_AWLEN   (hps_0_h2f_axi_master_awlen),   //               .awlen
		.h2f_AWSIZE  (hps_0_h2f_axi_master_awsize),  //               .awsize
		.h2f_AWBURST (hps_0_h2f_axi_master_awburst), //               .awburst
		.h2f_AWLOCK  (hps_0_h2f_axi_master_awlock),  //               .awlock
		.h2f_AWCACHE (hps_0_h2f_axi_master_awcache), //               .awcache
		.h2f_AWPROT  (hps_0_h2f_axi_master_awprot),  //               .awprot
		.h2f_AWVALID (hps_0_h2f_axi_master_awvalid), //               .awvalid
		.h2f_AWREADY (hps_0_h2f_axi_master_awready), //               .awready
		.h2f_WID     (hps_0_h2f_axi_master_wid),     //               .wid
		.h2f_WDATA   (hps_0_h2f_axi_master_wdata),   //               .wdata
		.h2f_WSTRB   (hps_0_h2f_axi_master_wstrb),   //               .wstrb
		.h2f_WLAST   (hps_0_h2f_axi_master_wlast),   //               .wlast
		.h2f_WVALID  (hps_0_h2f_axi_master_wvalid),  //               .wvalid
		.h2f_WREADY  (hps_0_h2f_axi_master_wready),  //               .wready
		.h2f_BID     (hps_0_h2f_axi_master_bid),     //               .bid
		.h2f_BRESP   (hps_0_h2f_axi_master_bresp),   //               .bresp
		.h2f_BVALID  (hps_0_h2f_axi_master_bvalid),  //               .bvalid
		.h2f_BREADY  (hps_0_h2f_axi_master_bready),  //               .bready
		.h2f_ARID    (hps_0_h2f_axi_master_arid),    //               .arid
		.h2f_ARADDR  (hps_0_h2f_axi_master_araddr),  //               .araddr
		.h2f_ARLEN   (hps_0_h2f_axi_master_arlen),   //               .arlen
		.h2f_ARSIZE  (hps_0_h2f_axi_master_arsize),  //               .arsize
		.h2f_ARBURST (hps_0_h2f_axi_master_arburst), //               .arburst
		.h2f_ARLOCK  (hps_0_h2f_axi_master_arlock),  //               .arlock
		.h2f_ARCACHE (hps_0_h2f_axi_master_arcache), //               .arcache
		.h2f_ARPROT  (hps_0_h2f_axi_master_arprot),  //               .arprot
		.h2f_ARVALID (hps_0_h2f_axi_master_arvalid), //               .arvalid
		.h2f_ARREADY (hps_0_h2f_axi_master_arready), //               .arready
		.h2f_RID     (hps_0_h2f_axi_master_rid),     //               .rid
		.h2f_RDATA   (hps_0_h2f_axi_master_rdata),   //               .rdata
		.h2f_RRESP   (hps_0_h2f_axi_master_rresp),   //               .rresp
		.h2f_RLAST   (hps_0_h2f_axi_master_rlast),   //               .rlast
		.h2f_RVALID  (hps_0_h2f_axi_master_rvalid),  //               .rvalid
		.h2f_RREADY  (hps_0_h2f_axi_master_rready)   //               .rready
	);

	jaxa_autoStart linkdisable (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_linkdisable_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_linkdisable_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_linkdisable_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_linkdisable_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_linkdisable_s1_readdata),   //                    .readdata
		.out_port   (linkdisable_external_connection_export)       // external_connection.export
	);

	jaxa_autoStart linkstart (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_linkstart_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_linkstart_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_linkstart_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_linkstart_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_linkstart_s1_readdata),   //                    .readdata
		.out_port   (linkstart_external_connection_export)       // external_connection.export
	);

	jaxa_linkStatus linkstatus (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_linkstatus_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_linkstatus_s1_readdata), //                    .readdata
		.in_port  (linkstatus_external_connection_export)     // external_connection.export
	);

	jaxa_creditCount outstandingcount (
		.clk      (clk_clk),                                        //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address  (mm_interconnect_0_outstandingcount_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_outstandingcount_s1_readdata), //                    .readdata
		.in_port  (outstandingcount_external_connection_export)     // external_connection.export
	);

	jaxa_pll_0 pll_0 (
		.refclk   (clk_clk),                //  refclk.clk
		.rst      (~hps_0_h2f_reset_reset), //   reset.reset
		.outclk_0 (pll_0_outclk0_clk),      // outclk0.clk
		.locked   ()                        //  locked.export
	);

	jaxa_receiveActivity receiveactivity (
		.clk      (clk_clk),                                       //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address  (mm_interconnect_0_receiveactivity_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_receiveactivity_s1_readdata), //                    .readdata
		.in_port  (receiveactivity_external_connection_export)     // external_connection.export
	);

	jaxa_autoStart receiveclock (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_receiveclock_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_receiveclock_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_receiveclock_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_receiveclock_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_receiveclock_s1_readdata),   //                    .readdata
		.out_port   (receiveclock_external_connection_export)       // external_connection.export
	);

	jaxa_receiveActivity receivefifodatacount (
		.clk      (clk_clk),                                            //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                    //               reset.reset_n
		.address  (mm_interconnect_0_receivefifodatacount_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_receivefifodatacount_s1_readdata), //                    .readdata
		.in_port  (receivefifodatacount_external_connection_export)     // external_connection.export
	);

	jaxa_receiveFIFODataOut receivefifodataout (
		.clk      (clk_clk),                                          //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address  (mm_interconnect_0_receivefifodataout_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_receivefifodataout_s1_readdata), //                    .readdata
		.in_port  (receivefifodataout_external_connection_export)     // external_connection.export
	);

	jaxa_receiveActivity receivefifoempty (
		.clk      (clk_clk),                                        //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address  (mm_interconnect_0_receivefifoempty_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_receivefifoempty_s1_readdata), //                    .readdata
		.in_port  (receivefifoempty_external_connection_export)     // external_connection.export
	);

	jaxa_receiveActivity receivefifofull (
		.clk      (clk_clk),                                       //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address  (mm_interconnect_0_receivefifofull_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_receivefifofull_s1_readdata), //                    .readdata
		.in_port  (receivefifofull_external_connection_export)     // external_connection.export
	);

	jaxa_autoStart receivefiforeadenable (
		.clk        (clk_clk),                                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                       //               reset.reset_n
		.address    (mm_interconnect_0_receivefiforeadenable_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_receivefiforeadenable_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_receivefiforeadenable_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_receivefiforeadenable_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_receivefiforeadenable_s1_readdata),   //                    .readdata
		.out_port   (receivefiforeadenable_external_connection_export)       // external_connection.export
	);

	jaxa_autoStart spacewiredatain (
		.clk        (clk_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_spacewiredatain_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_spacewiredatain_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_spacewiredatain_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_spacewiredatain_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_spacewiredatain_s1_readdata),   //                    .readdata
		.out_port   (spacewiredatain_external_connection_export)       // external_connection.export
	);

	jaxa_receiveActivity spacewiredataout (
		.clk      (clk_clk),                                        //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address  (mm_interconnect_0_spacewiredataout_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_spacewiredataout_s1_readdata), //                    .readdata
		.in_port  (spacewiredataout_external_connection_export)     // external_connection.export
	);

	jaxa_autoStart spacewirestrobein (
		.clk        (clk_clk),                                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (mm_interconnect_0_spacewirestrobein_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_spacewirestrobein_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_spacewirestrobein_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_spacewirestrobein_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_spacewirestrobein_s1_readdata),   //                    .readdata
		.out_port   (spacewirestrobein_external_connection_export)       // external_connection.export
	);

	jaxa_receiveActivity spacewirestrobeout (
		.clk      (clk_clk),                                          //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address  (mm_interconnect_0_spacewirestrobeout_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_spacewirestrobeout_s1_readdata), //                    .readdata
		.in_port  (spacewirestrobeout_external_connection_export)     // external_connection.export
	);

	jaxa_autoStart statisticalinformationclear (
		.clk        (clk_clk),                                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                             //               reset.reset_n
		.address    (mm_interconnect_0_statisticalinformationclear_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_statisticalinformationclear_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_statisticalinformationclear_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_statisticalinformationclear_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_statisticalinformationclear_s1_readdata),   //                    .readdata
		.out_port   (statisticalinformationclear_external_connection_export)       // external_connection.export
	);

	jaxa_statisticalInformation_0 statisticalinformation_0 (
		.clk      (clk_clk),                                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                        //               reset.reset_n
		.address  (mm_interconnect_0_statisticalinformation_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_statisticalinformation_0_s1_readdata), //                    .readdata
		.in_port  (statisticalinformation_0_external_connection_export)     // external_connection.export
	);

	jaxa_statisticalInformation_1 statisticalinformation_1 (
		.clk        (clk_clk),                                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                          //               reset.reset_n
		.address    (mm_interconnect_0_statisticalinformation_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_statisticalinformation_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_statisticalinformation_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_statisticalinformation_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_statisticalinformation_1_s1_readdata),   //                    .readdata
		.out_port   (statisticalinformation_1_external_connection_export)       // external_connection.export
	);

	jaxa_autoStart tickin (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_tickin_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_tickin_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_tickin_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_tickin_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_tickin_s1_readdata),   //                    .readdata
		.out_port   (tickin_external_connection_export)       // external_connection.export
	);

	jaxa_receiveActivity tickout (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_tickout_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_tickout_s1_readdata), //                    .readdata
		.in_port  (tickout_external_connection_export)     // external_connection.export
	);

	jaxa_timeIn timein (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_timein_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_timein_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_timein_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_timein_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_timein_s1_readdata),   //                    .readdata
		.out_port   (timein_external_connection_export)       // external_connection.export
	);

	jaxa_creditCount timeout (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_timeout_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_timeout_s1_readdata), //                    .readdata
		.in_port  (timeout_external_connection_export)     // external_connection.export
	);

	jaxa_receiveActivity transmitactivity (
		.clk      (clk_clk),                                        //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address  (mm_interconnect_0_transmitactivity_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_transmitactivity_s1_readdata), //                    .readdata
		.in_port  (transmitactivity_external_connection_export)     // external_connection.export
	);

	jaxa_autoStart transmitclock (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_transmitclock_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_transmitclock_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_transmitclock_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_transmitclock_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_transmitclock_s1_readdata),   //                    .readdata
		.out_port   (transmitclock_external_connection_export)       // external_connection.export
	);

	jaxa_timeIn transmitclockdividevalue (
		.clk        (clk_clk),                                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                          //               reset.reset_n
		.address    (mm_interconnect_0_transmitclockdividevalue_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_transmitclockdividevalue_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_transmitclockdividevalue_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_transmitclockdividevalue_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_transmitclockdividevalue_s1_readdata),   //                    .readdata
		.out_port   (transmitclockdividevalue_external_connection_export)       // external_connection.export
	);

	jaxa_creditCount transmitfifodatacount (
		.clk      (clk_clk),                                             //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                     //               reset.reset_n
		.address  (mm_interconnect_0_transmitfifodatacount_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_transmitfifodatacount_s1_readdata), //                    .readdata
		.in_port  (transmitfifodatacount_external_connection_export)     // external_connection.export
	);

	jaxa_transmitFIFODataIn transmitfifodatain (
		.clk        (clk_clk),                                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                    //               reset.reset_n
		.address    (mm_interconnect_0_transmitfifodatain_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_transmitfifodatain_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_transmitfifodatain_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_transmitfifodatain_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_transmitfifodatain_s1_readdata),   //                    .readdata
		.out_port   (transmitfifodatain_external_connection_export)       // external_connection.export
	);

	jaxa_receiveActivity transmitfifofull (
		.clk      (clk_clk),                                        //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address  (mm_interconnect_0_transmitfifofull_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_transmitfifofull_s1_readdata), //                    .readdata
		.in_port  (transmitfifofull_external_connection_export)     // external_connection.export
	);

	jaxa_autoStart transmitfifowriteenable (
		.clk        (clk_clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                         //               reset.reset_n
		.address    (mm_interconnect_0_transmitfifowriteenable_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_transmitfifowriteenable_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_transmitfifowriteenable_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_transmitfifowriteenable_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_transmitfifowriteenable_s1_readdata),   //                    .readdata
		.out_port   (transmitfifowriteenable_external_connection_export)       // external_connection.export
	);

	jaxa_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_h2f_axi_master_awid                                        (hps_0_h2f_axi_master_awid),                                   //                                       hps_0_h2f_axi_master.awid
		.hps_0_h2f_axi_master_awaddr                                      (hps_0_h2f_axi_master_awaddr),                                 //                                                           .awaddr
		.hps_0_h2f_axi_master_awlen                                       (hps_0_h2f_axi_master_awlen),                                  //                                                           .awlen
		.hps_0_h2f_axi_master_awsize                                      (hps_0_h2f_axi_master_awsize),                                 //                                                           .awsize
		.hps_0_h2f_axi_master_awburst                                     (hps_0_h2f_axi_master_awburst),                                //                                                           .awburst
		.hps_0_h2f_axi_master_awlock                                      (hps_0_h2f_axi_master_awlock),                                 //                                                           .awlock
		.hps_0_h2f_axi_master_awcache                                     (hps_0_h2f_axi_master_awcache),                                //                                                           .awcache
		.hps_0_h2f_axi_master_awprot                                      (hps_0_h2f_axi_master_awprot),                                 //                                                           .awprot
		.hps_0_h2f_axi_master_awvalid                                     (hps_0_h2f_axi_master_awvalid),                                //                                                           .awvalid
		.hps_0_h2f_axi_master_awready                                     (hps_0_h2f_axi_master_awready),                                //                                                           .awready
		.hps_0_h2f_axi_master_wid                                         (hps_0_h2f_axi_master_wid),                                    //                                                           .wid
		.hps_0_h2f_axi_master_wdata                                       (hps_0_h2f_axi_master_wdata),                                  //                                                           .wdata
		.hps_0_h2f_axi_master_wstrb                                       (hps_0_h2f_axi_master_wstrb),                                  //                                                           .wstrb
		.hps_0_h2f_axi_master_wlast                                       (hps_0_h2f_axi_master_wlast),                                  //                                                           .wlast
		.hps_0_h2f_axi_master_wvalid                                      (hps_0_h2f_axi_master_wvalid),                                 //                                                           .wvalid
		.hps_0_h2f_axi_master_wready                                      (hps_0_h2f_axi_master_wready),                                 //                                                           .wready
		.hps_0_h2f_axi_master_bid                                         (hps_0_h2f_axi_master_bid),                                    //                                                           .bid
		.hps_0_h2f_axi_master_bresp                                       (hps_0_h2f_axi_master_bresp),                                  //                                                           .bresp
		.hps_0_h2f_axi_master_bvalid                                      (hps_0_h2f_axi_master_bvalid),                                 //                                                           .bvalid
		.hps_0_h2f_axi_master_bready                                      (hps_0_h2f_axi_master_bready),                                 //                                                           .bready
		.hps_0_h2f_axi_master_arid                                        (hps_0_h2f_axi_master_arid),                                   //                                                           .arid
		.hps_0_h2f_axi_master_araddr                                      (hps_0_h2f_axi_master_araddr),                                 //                                                           .araddr
		.hps_0_h2f_axi_master_arlen                                       (hps_0_h2f_axi_master_arlen),                                  //                                                           .arlen
		.hps_0_h2f_axi_master_arsize                                      (hps_0_h2f_axi_master_arsize),                                 //                                                           .arsize
		.hps_0_h2f_axi_master_arburst                                     (hps_0_h2f_axi_master_arburst),                                //                                                           .arburst
		.hps_0_h2f_axi_master_arlock                                      (hps_0_h2f_axi_master_arlock),                                 //                                                           .arlock
		.hps_0_h2f_axi_master_arcache                                     (hps_0_h2f_axi_master_arcache),                                //                                                           .arcache
		.hps_0_h2f_axi_master_arprot                                      (hps_0_h2f_axi_master_arprot),                                 //                                                           .arprot
		.hps_0_h2f_axi_master_arvalid                                     (hps_0_h2f_axi_master_arvalid),                                //                                                           .arvalid
		.hps_0_h2f_axi_master_arready                                     (hps_0_h2f_axi_master_arready),                                //                                                           .arready
		.hps_0_h2f_axi_master_rid                                         (hps_0_h2f_axi_master_rid),                                    //                                                           .rid
		.hps_0_h2f_axi_master_rdata                                       (hps_0_h2f_axi_master_rdata),                                  //                                                           .rdata
		.hps_0_h2f_axi_master_rresp                                       (hps_0_h2f_axi_master_rresp),                                  //                                                           .rresp
		.hps_0_h2f_axi_master_rlast                                       (hps_0_h2f_axi_master_rlast),                                  //                                                           .rlast
		.hps_0_h2f_axi_master_rvalid                                      (hps_0_h2f_axi_master_rvalid),                                 //                                                           .rvalid
		.hps_0_h2f_axi_master_rready                                      (hps_0_h2f_axi_master_rready),                                 //                                                           .rready
		.clk_0_clk_clk                                                    (clk_clk),                                                     //                                                  clk_0_clk.clk
		.autoStart_reset_reset_bridge_in_reset_reset                      (rst_controller_reset_out_reset),                              //                      autoStart_reset_reset_bridge_in_reset.reset
		.hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                          // hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.autoStart_s1_address                                             (mm_interconnect_0_autostart_s1_address),                      //                                               autoStart_s1.address
		.autoStart_s1_write                                               (mm_interconnect_0_autostart_s1_write),                        //                                                           .write
		.autoStart_s1_readdata                                            (mm_interconnect_0_autostart_s1_readdata),                     //                                                           .readdata
		.autoStart_s1_writedata                                           (mm_interconnect_0_autostart_s1_writedata),                    //                                                           .writedata
		.autoStart_s1_chipselect                                          (mm_interconnect_0_autostart_s1_chipselect),                   //                                                           .chipselect
		.controlFlagsIn_s1_address                                        (mm_interconnect_0_controlflagsin_s1_address),                 //                                          controlFlagsIn_s1.address
		.controlFlagsIn_s1_write                                          (mm_interconnect_0_controlflagsin_s1_write),                   //                                                           .write
		.controlFlagsIn_s1_readdata                                       (mm_interconnect_0_controlflagsin_s1_readdata),                //                                                           .readdata
		.controlFlagsIn_s1_writedata                                      (mm_interconnect_0_controlflagsin_s1_writedata),               //                                                           .writedata
		.controlFlagsIn_s1_chipselect                                     (mm_interconnect_0_controlflagsin_s1_chipselect),              //                                                           .chipselect
		.controlFlagsOut_s1_address                                       (mm_interconnect_0_controlflagsout_s1_address),                //                                         controlFlagsOut_s1.address
		.controlFlagsOut_s1_readdata                                      (mm_interconnect_0_controlflagsout_s1_readdata),               //                                                           .readdata
		.creditCount_s1_address                                           (mm_interconnect_0_creditcount_s1_address),                    //                                             creditCount_s1.address
		.creditCount_s1_readdata                                          (mm_interconnect_0_creditcount_s1_readdata),                   //                                                           .readdata
		.errorStatus_s1_address                                           (mm_interconnect_0_errorstatus_s1_address),                    //                                             errorStatus_s1.address
		.errorStatus_s1_readdata                                          (mm_interconnect_0_errorstatus_s1_readdata),                   //                                                           .readdata
		.linkDisable_s1_address                                           (mm_interconnect_0_linkdisable_s1_address),                    //                                             linkDisable_s1.address
		.linkDisable_s1_write                                             (mm_interconnect_0_linkdisable_s1_write),                      //                                                           .write
		.linkDisable_s1_readdata                                          (mm_interconnect_0_linkdisable_s1_readdata),                   //                                                           .readdata
		.linkDisable_s1_writedata                                         (mm_interconnect_0_linkdisable_s1_writedata),                  //                                                           .writedata
		.linkDisable_s1_chipselect                                        (mm_interconnect_0_linkdisable_s1_chipselect),                 //                                                           .chipselect
		.linkStart_s1_address                                             (mm_interconnect_0_linkstart_s1_address),                      //                                               linkStart_s1.address
		.linkStart_s1_write                                               (mm_interconnect_0_linkstart_s1_write),                        //                                                           .write
		.linkStart_s1_readdata                                            (mm_interconnect_0_linkstart_s1_readdata),                     //                                                           .readdata
		.linkStart_s1_writedata                                           (mm_interconnect_0_linkstart_s1_writedata),                    //                                                           .writedata
		.linkStart_s1_chipselect                                          (mm_interconnect_0_linkstart_s1_chipselect),                   //                                                           .chipselect
		.linkStatus_s1_address                                            (mm_interconnect_0_linkstatus_s1_address),                     //                                              linkStatus_s1.address
		.linkStatus_s1_readdata                                           (mm_interconnect_0_linkstatus_s1_readdata),                    //                                                           .readdata
		.outstandingCount_s1_address                                      (mm_interconnect_0_outstandingcount_s1_address),               //                                        outstandingCount_s1.address
		.outstandingCount_s1_readdata                                     (mm_interconnect_0_outstandingcount_s1_readdata),              //                                                           .readdata
		.receiveActivity_s1_address                                       (mm_interconnect_0_receiveactivity_s1_address),                //                                         receiveActivity_s1.address
		.receiveActivity_s1_readdata                                      (mm_interconnect_0_receiveactivity_s1_readdata),               //                                                           .readdata
		.receiveClock_s1_address                                          (mm_interconnect_0_receiveclock_s1_address),                   //                                            receiveClock_s1.address
		.receiveClock_s1_write                                            (mm_interconnect_0_receiveclock_s1_write),                     //                                                           .write
		.receiveClock_s1_readdata                                         (mm_interconnect_0_receiveclock_s1_readdata),                  //                                                           .readdata
		.receiveClock_s1_writedata                                        (mm_interconnect_0_receiveclock_s1_writedata),                 //                                                           .writedata
		.receiveClock_s1_chipselect                                       (mm_interconnect_0_receiveclock_s1_chipselect),                //                                                           .chipselect
		.receiveFIFODataCount_s1_address                                  (mm_interconnect_0_receivefifodatacount_s1_address),           //                                    receiveFIFODataCount_s1.address
		.receiveFIFODataCount_s1_readdata                                 (mm_interconnect_0_receivefifodatacount_s1_readdata),          //                                                           .readdata
		.receiveFIFODataOut_s1_address                                    (mm_interconnect_0_receivefifodataout_s1_address),             //                                      receiveFIFODataOut_s1.address
		.receiveFIFODataOut_s1_readdata                                   (mm_interconnect_0_receivefifodataout_s1_readdata),            //                                                           .readdata
		.receiveFIFOEmpty_s1_address                                      (mm_interconnect_0_receivefifoempty_s1_address),               //                                        receiveFIFOEmpty_s1.address
		.receiveFIFOEmpty_s1_readdata                                     (mm_interconnect_0_receivefifoempty_s1_readdata),              //                                                           .readdata
		.receiveFIFOFull_s1_address                                       (mm_interconnect_0_receivefifofull_s1_address),                //                                         receiveFIFOFull_s1.address
		.receiveFIFOFull_s1_readdata                                      (mm_interconnect_0_receivefifofull_s1_readdata),               //                                                           .readdata
		.receiveFIFOReadEnable_s1_address                                 (mm_interconnect_0_receivefiforeadenable_s1_address),          //                                   receiveFIFOReadEnable_s1.address
		.receiveFIFOReadEnable_s1_write                                   (mm_interconnect_0_receivefiforeadenable_s1_write),            //                                                           .write
		.receiveFIFOReadEnable_s1_readdata                                (mm_interconnect_0_receivefiforeadenable_s1_readdata),         //                                                           .readdata
		.receiveFIFOReadEnable_s1_writedata                               (mm_interconnect_0_receivefiforeadenable_s1_writedata),        //                                                           .writedata
		.receiveFIFOReadEnable_s1_chipselect                              (mm_interconnect_0_receivefiforeadenable_s1_chipselect),       //                                                           .chipselect
		.spaceWireDataIn_s1_address                                       (mm_interconnect_0_spacewiredatain_s1_address),                //                                         spaceWireDataIn_s1.address
		.spaceWireDataIn_s1_write                                         (mm_interconnect_0_spacewiredatain_s1_write),                  //                                                           .write
		.spaceWireDataIn_s1_readdata                                      (mm_interconnect_0_spacewiredatain_s1_readdata),               //                                                           .readdata
		.spaceWireDataIn_s1_writedata                                     (mm_interconnect_0_spacewiredatain_s1_writedata),              //                                                           .writedata
		.spaceWireDataIn_s1_chipselect                                    (mm_interconnect_0_spacewiredatain_s1_chipselect),             //                                                           .chipselect
		.spaceWireDataOut_s1_address                                      (mm_interconnect_0_spacewiredataout_s1_address),               //                                        spaceWireDataOut_s1.address
		.spaceWireDataOut_s1_readdata                                     (mm_interconnect_0_spacewiredataout_s1_readdata),              //                                                           .readdata
		.spaceWireStrobeIn_s1_address                                     (mm_interconnect_0_spacewirestrobein_s1_address),              //                                       spaceWireStrobeIn_s1.address
		.spaceWireStrobeIn_s1_write                                       (mm_interconnect_0_spacewirestrobein_s1_write),                //                                                           .write
		.spaceWireStrobeIn_s1_readdata                                    (mm_interconnect_0_spacewirestrobein_s1_readdata),             //                                                           .readdata
		.spaceWireStrobeIn_s1_writedata                                   (mm_interconnect_0_spacewirestrobein_s1_writedata),            //                                                           .writedata
		.spaceWireStrobeIn_s1_chipselect                                  (mm_interconnect_0_spacewirestrobein_s1_chipselect),           //                                                           .chipselect
		.spaceWireStrobeOut_s1_address                                    (mm_interconnect_0_spacewirestrobeout_s1_address),             //                                      spaceWireStrobeOut_s1.address
		.spaceWireStrobeOut_s1_readdata                                   (mm_interconnect_0_spacewirestrobeout_s1_readdata),            //                                                           .readdata
		.statisticalInformation_0_s1_address                              (mm_interconnect_0_statisticalinformation_0_s1_address),       //                                statisticalInformation_0_s1.address
		.statisticalInformation_0_s1_readdata                             (mm_interconnect_0_statisticalinformation_0_s1_readdata),      //                                                           .readdata
		.statisticalInformation_1_s1_address                              (mm_interconnect_0_statisticalinformation_1_s1_address),       //                                statisticalInformation_1_s1.address
		.statisticalInformation_1_s1_write                                (mm_interconnect_0_statisticalinformation_1_s1_write),         //                                                           .write
		.statisticalInformation_1_s1_readdata                             (mm_interconnect_0_statisticalinformation_1_s1_readdata),      //                                                           .readdata
		.statisticalInformation_1_s1_writedata                            (mm_interconnect_0_statisticalinformation_1_s1_writedata),     //                                                           .writedata
		.statisticalInformation_1_s1_chipselect                           (mm_interconnect_0_statisticalinformation_1_s1_chipselect),    //                                                           .chipselect
		.statisticalInformationClear_s1_address                           (mm_interconnect_0_statisticalinformationclear_s1_address),    //                             statisticalInformationClear_s1.address
		.statisticalInformationClear_s1_write                             (mm_interconnect_0_statisticalinformationclear_s1_write),      //                                                           .write
		.statisticalInformationClear_s1_readdata                          (mm_interconnect_0_statisticalinformationclear_s1_readdata),   //                                                           .readdata
		.statisticalInformationClear_s1_writedata                         (mm_interconnect_0_statisticalinformationclear_s1_writedata),  //                                                           .writedata
		.statisticalInformationClear_s1_chipselect                        (mm_interconnect_0_statisticalinformationclear_s1_chipselect), //                                                           .chipselect
		.tickIn_s1_address                                                (mm_interconnect_0_tickin_s1_address),                         //                                                  tickIn_s1.address
		.tickIn_s1_write                                                  (mm_interconnect_0_tickin_s1_write),                           //                                                           .write
		.tickIn_s1_readdata                                               (mm_interconnect_0_tickin_s1_readdata),                        //                                                           .readdata
		.tickIn_s1_writedata                                              (mm_interconnect_0_tickin_s1_writedata),                       //                                                           .writedata
		.tickIn_s1_chipselect                                             (mm_interconnect_0_tickin_s1_chipselect),                      //                                                           .chipselect
		.tickOut_s1_address                                               (mm_interconnect_0_tickout_s1_address),                        //                                                 tickOut_s1.address
		.tickOut_s1_readdata                                              (mm_interconnect_0_tickout_s1_readdata),                       //                                                           .readdata
		.timeIn_s1_address                                                (mm_interconnect_0_timein_s1_address),                         //                                                  timeIn_s1.address
		.timeIn_s1_write                                                  (mm_interconnect_0_timein_s1_write),                           //                                                           .write
		.timeIn_s1_readdata                                               (mm_interconnect_0_timein_s1_readdata),                        //                                                           .readdata
		.timeIn_s1_writedata                                              (mm_interconnect_0_timein_s1_writedata),                       //                                                           .writedata
		.timeIn_s1_chipselect                                             (mm_interconnect_0_timein_s1_chipselect),                      //                                                           .chipselect
		.timeOut_s1_address                                               (mm_interconnect_0_timeout_s1_address),                        //                                                 timeOut_s1.address
		.timeOut_s1_readdata                                              (mm_interconnect_0_timeout_s1_readdata),                       //                                                           .readdata
		.transmitActivity_s1_address                                      (mm_interconnect_0_transmitactivity_s1_address),               //                                        transmitActivity_s1.address
		.transmitActivity_s1_readdata                                     (mm_interconnect_0_transmitactivity_s1_readdata),              //                                                           .readdata
		.transmitClock_s1_address                                         (mm_interconnect_0_transmitclock_s1_address),                  //                                           transmitClock_s1.address
		.transmitClock_s1_write                                           (mm_interconnect_0_transmitclock_s1_write),                    //                                                           .write
		.transmitClock_s1_readdata                                        (mm_interconnect_0_transmitclock_s1_readdata),                 //                                                           .readdata
		.transmitClock_s1_writedata                                       (mm_interconnect_0_transmitclock_s1_writedata),                //                                                           .writedata
		.transmitClock_s1_chipselect                                      (mm_interconnect_0_transmitclock_s1_chipselect),               //                                                           .chipselect
		.transmitClockDivideValue_s1_address                              (mm_interconnect_0_transmitclockdividevalue_s1_address),       //                                transmitClockDivideValue_s1.address
		.transmitClockDivideValue_s1_write                                (mm_interconnect_0_transmitclockdividevalue_s1_write),         //                                                           .write
		.transmitClockDivideValue_s1_readdata                             (mm_interconnect_0_transmitclockdividevalue_s1_readdata),      //                                                           .readdata
		.transmitClockDivideValue_s1_writedata                            (mm_interconnect_0_transmitclockdividevalue_s1_writedata),     //                                                           .writedata
		.transmitClockDivideValue_s1_chipselect                           (mm_interconnect_0_transmitclockdividevalue_s1_chipselect),    //                                                           .chipselect
		.transmitFIFODataCount_s1_address                                 (mm_interconnect_0_transmitfifodatacount_s1_address),          //                                   transmitFIFODataCount_s1.address
		.transmitFIFODataCount_s1_readdata                                (mm_interconnect_0_transmitfifodatacount_s1_readdata),         //                                                           .readdata
		.transmitFIFODataIn_s1_address                                    (mm_interconnect_0_transmitfifodatain_s1_address),             //                                      transmitFIFODataIn_s1.address
		.transmitFIFODataIn_s1_write                                      (mm_interconnect_0_transmitfifodatain_s1_write),               //                                                           .write
		.transmitFIFODataIn_s1_readdata                                   (mm_interconnect_0_transmitfifodatain_s1_readdata),            //                                                           .readdata
		.transmitFIFODataIn_s1_writedata                                  (mm_interconnect_0_transmitfifodatain_s1_writedata),           //                                                           .writedata
		.transmitFIFODataIn_s1_chipselect                                 (mm_interconnect_0_transmitfifodatain_s1_chipselect),          //                                                           .chipselect
		.transmitFIFOFull_s1_address                                      (mm_interconnect_0_transmitfifofull_s1_address),               //                                        transmitFIFOFull_s1.address
		.transmitFIFOFull_s1_readdata                                     (mm_interconnect_0_transmitfifofull_s1_readdata),              //                                                           .readdata
		.transmitFIFOWriteEnable_s1_address                               (mm_interconnect_0_transmitfifowriteenable_s1_address),        //                                 transmitFIFOWriteEnable_s1.address
		.transmitFIFOWriteEnable_s1_write                                 (mm_interconnect_0_transmitfifowriteenable_s1_write),          //                                                           .write
		.transmitFIFOWriteEnable_s1_readdata                              (mm_interconnect_0_transmitfifowriteenable_s1_readdata),       //                                                           .readdata
		.transmitFIFOWriteEnable_s1_writedata                             (mm_interconnect_0_transmitfifowriteenable_s1_writedata),      //                                                           .writedata
		.transmitFIFOWriteEnable_s1_chipselect                            (mm_interconnect_0_transmitfifowriteenable_s1_chipselect)      //                                                           .chipselect
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~hps_0_h2f_reset_reset),         // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~hps_0_h2f_reset_reset),             // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
