// spw_light.v

// Generated using ACDS version 17.1 593

`timescale 1 ps / 1 ps
module spw_light (
		output wire        autostart_external_connection_export,  //  autostart_external_connection.export
		input  wire        clk_clk,                               //                            clk.clk
		input  wire        connecting_external_connection_export, // connecting_external_connection.export
		output wire [1:0]  ctrl_in_external_connection_export,    //    ctrl_in_external_connection.export
		input  wire [1:0]  ctrl_out_external_connection_export,   //   ctrl_out_external_connection.export
		input  wire        errcred_external_connection_export,    //    errcred_external_connection.export
		input  wire        errdisc_external_connection_export,    //    errdisc_external_connection.export
		input  wire        erresc_external_connection_export,     //     erresc_external_connection.export
		input  wire        errpar_external_connection_export,     //     errpar_external_connection.export
		output wire        linkdis_external_connection_export,    //    linkdis_external_connection.export
		output wire        linkstart_external_connection_export,  //  linkstart_external_connection.export
		output wire [12:0] memory_mem_a,                          //                         memory.mem_a
		output wire [2:0]  memory_mem_ba,                         //                               .mem_ba
		output wire        memory_mem_ck,                         //                               .mem_ck
		output wire        memory_mem_ck_n,                       //                               .mem_ck_n
		output wire        memory_mem_cke,                        //                               .mem_cke
		output wire        memory_mem_cs_n,                       //                               .mem_cs_n
		output wire        memory_mem_ras_n,                      //                               .mem_ras_n
		output wire        memory_mem_cas_n,                      //                               .mem_cas_n
		output wire        memory_mem_we_n,                       //                               .mem_we_n
		output wire        memory_mem_reset_n,                    //                               .mem_reset_n
		inout  wire [7:0]  memory_mem_dq,                         //                               .mem_dq
		inout  wire        memory_mem_dqs,                        //                               .mem_dqs
		inout  wire        memory_mem_dqs_n,                      //                               .mem_dqs_n
		output wire        memory_mem_odt,                        //                               .mem_odt
		output wire        memory_mem_dm,                         //                               .mem_dm
		input  wire        memory_oct_rzqin,                      //                               .oct_rzqin
		output wire        pll_0_locked_export,                   //                   pll_0_locked.export
		output wire        pll_0_outclk0_clk,                     //                  pll_0_outclk0.clk
		input  wire        reset_reset_n,                         //                          reset.reset_n
		input  wire        running_external_connection_export,    //    running_external_connection.export
		input  wire [7:0]  rxdata_external_connection_export,     //     rxdata_external_connection.export
		input  wire        rxflag_external_connection_export,     //     rxflag_external_connection.export
		input  wire        rxhalff_external_connection_export,    //    rxhalff_external_connection.export
		output wire        rxread_external_connection_export,     //     rxread_external_connection.export
		input  wire        rxvalid_external_connection_export,    //    rxvalid_external_connection.export
		input  wire        started_external_connection_export,    //    started_external_connection.export
		output wire        tick_in_external_connection_export,    //    tick_in_external_connection.export
		input  wire        tick_out_external_connection_export,   //   tick_out_external_connection.export
		output wire [5:0]  time_in_external_connection_export,    //    time_in_external_connection.export
		input  wire [5:0]  time_out_external_connection_export,   //   time_out_external_connection.export
		output wire [7:0]  txdata_external_connection_export,     //     txdata_external_connection.export
		output wire [7:0]  txdivcnt_external_connection_export,   //   txdivcnt_external_connection.export
		output wire        txflag_external_connection_export,     //     txflag_external_connection.export
		input  wire        txhalff_external_connection_export,    //    txhalff_external_connection.export
		input  wire        txrdy_external_connection_export,      //      txrdy_external_connection.export
		output wire        txwrite_external_connection_export     //    txwrite_external_connection.export
	);

	wire   [1:0] hps_0_h2f_axi_master_awburst;              // hps_0:h2f_AWBURST -> mm_interconnect_0:hps_0_h2f_axi_master_awburst
	wire   [3:0] hps_0_h2f_axi_master_arlen;                // hps_0:h2f_ARLEN -> mm_interconnect_0:hps_0_h2f_axi_master_arlen
	wire   [3:0] hps_0_h2f_axi_master_wstrb;                // hps_0:h2f_WSTRB -> mm_interconnect_0:hps_0_h2f_axi_master_wstrb
	wire         hps_0_h2f_axi_master_wready;               // mm_interconnect_0:hps_0_h2f_axi_master_wready -> hps_0:h2f_WREADY
	wire  [11:0] hps_0_h2f_axi_master_rid;                  // mm_interconnect_0:hps_0_h2f_axi_master_rid -> hps_0:h2f_RID
	wire         hps_0_h2f_axi_master_rready;               // hps_0:h2f_RREADY -> mm_interconnect_0:hps_0_h2f_axi_master_rready
	wire   [3:0] hps_0_h2f_axi_master_awlen;                // hps_0:h2f_AWLEN -> mm_interconnect_0:hps_0_h2f_axi_master_awlen
	wire  [11:0] hps_0_h2f_axi_master_wid;                  // hps_0:h2f_WID -> mm_interconnect_0:hps_0_h2f_axi_master_wid
	wire   [3:0] hps_0_h2f_axi_master_arcache;              // hps_0:h2f_ARCACHE -> mm_interconnect_0:hps_0_h2f_axi_master_arcache
	wire         hps_0_h2f_axi_master_wvalid;               // hps_0:h2f_WVALID -> mm_interconnect_0:hps_0_h2f_axi_master_wvalid
	wire  [29:0] hps_0_h2f_axi_master_araddr;               // hps_0:h2f_ARADDR -> mm_interconnect_0:hps_0_h2f_axi_master_araddr
	wire   [2:0] hps_0_h2f_axi_master_arprot;               // hps_0:h2f_ARPROT -> mm_interconnect_0:hps_0_h2f_axi_master_arprot
	wire   [2:0] hps_0_h2f_axi_master_awprot;               // hps_0:h2f_AWPROT -> mm_interconnect_0:hps_0_h2f_axi_master_awprot
	wire  [31:0] hps_0_h2f_axi_master_wdata;                // hps_0:h2f_WDATA -> mm_interconnect_0:hps_0_h2f_axi_master_wdata
	wire         hps_0_h2f_axi_master_arvalid;              // hps_0:h2f_ARVALID -> mm_interconnect_0:hps_0_h2f_axi_master_arvalid
	wire   [3:0] hps_0_h2f_axi_master_awcache;              // hps_0:h2f_AWCACHE -> mm_interconnect_0:hps_0_h2f_axi_master_awcache
	wire  [11:0] hps_0_h2f_axi_master_arid;                 // hps_0:h2f_ARID -> mm_interconnect_0:hps_0_h2f_axi_master_arid
	wire   [1:0] hps_0_h2f_axi_master_arlock;               // hps_0:h2f_ARLOCK -> mm_interconnect_0:hps_0_h2f_axi_master_arlock
	wire   [1:0] hps_0_h2f_axi_master_awlock;               // hps_0:h2f_AWLOCK -> mm_interconnect_0:hps_0_h2f_axi_master_awlock
	wire  [29:0] hps_0_h2f_axi_master_awaddr;               // hps_0:h2f_AWADDR -> mm_interconnect_0:hps_0_h2f_axi_master_awaddr
	wire   [1:0] hps_0_h2f_axi_master_bresp;                // mm_interconnect_0:hps_0_h2f_axi_master_bresp -> hps_0:h2f_BRESP
	wire         hps_0_h2f_axi_master_arready;              // mm_interconnect_0:hps_0_h2f_axi_master_arready -> hps_0:h2f_ARREADY
	wire  [31:0] hps_0_h2f_axi_master_rdata;                // mm_interconnect_0:hps_0_h2f_axi_master_rdata -> hps_0:h2f_RDATA
	wire         hps_0_h2f_axi_master_awready;              // mm_interconnect_0:hps_0_h2f_axi_master_awready -> hps_0:h2f_AWREADY
	wire   [1:0] hps_0_h2f_axi_master_arburst;              // hps_0:h2f_ARBURST -> mm_interconnect_0:hps_0_h2f_axi_master_arburst
	wire   [2:0] hps_0_h2f_axi_master_arsize;               // hps_0:h2f_ARSIZE -> mm_interconnect_0:hps_0_h2f_axi_master_arsize
	wire         hps_0_h2f_axi_master_bready;               // hps_0:h2f_BREADY -> mm_interconnect_0:hps_0_h2f_axi_master_bready
	wire         hps_0_h2f_axi_master_rlast;                // mm_interconnect_0:hps_0_h2f_axi_master_rlast -> hps_0:h2f_RLAST
	wire         hps_0_h2f_axi_master_wlast;                // hps_0:h2f_WLAST -> mm_interconnect_0:hps_0_h2f_axi_master_wlast
	wire   [1:0] hps_0_h2f_axi_master_rresp;                // mm_interconnect_0:hps_0_h2f_axi_master_rresp -> hps_0:h2f_RRESP
	wire  [11:0] hps_0_h2f_axi_master_awid;                 // hps_0:h2f_AWID -> mm_interconnect_0:hps_0_h2f_axi_master_awid
	wire  [11:0] hps_0_h2f_axi_master_bid;                  // mm_interconnect_0:hps_0_h2f_axi_master_bid -> hps_0:h2f_BID
	wire         hps_0_h2f_axi_master_bvalid;               // mm_interconnect_0:hps_0_h2f_axi_master_bvalid -> hps_0:h2f_BVALID
	wire   [2:0] hps_0_h2f_axi_master_awsize;               // hps_0:h2f_AWSIZE -> mm_interconnect_0:hps_0_h2f_axi_master_awsize
	wire         hps_0_h2f_axi_master_awvalid;              // hps_0:h2f_AWVALID -> mm_interconnect_0:hps_0_h2f_axi_master_awvalid
	wire         hps_0_h2f_axi_master_rvalid;               // mm_interconnect_0:hps_0_h2f_axi_master_rvalid -> hps_0:h2f_RVALID
	wire         mm_interconnect_0_autostart_s1_chipselect; // mm_interconnect_0:autostart_s1_chipselect -> autostart:chipselect
	wire  [31:0] mm_interconnect_0_autostart_s1_readdata;   // autostart:readdata -> mm_interconnect_0:autostart_s1_readdata
	wire   [1:0] mm_interconnect_0_autostart_s1_address;    // mm_interconnect_0:autostart_s1_address -> autostart:address
	wire         mm_interconnect_0_autostart_s1_write;      // mm_interconnect_0:autostart_s1_write -> autostart:write_n
	wire  [31:0] mm_interconnect_0_autostart_s1_writedata;  // mm_interconnect_0:autostart_s1_writedata -> autostart:writedata
	wire         mm_interconnect_0_linkdis_s1_chipselect;   // mm_interconnect_0:linkdis_s1_chipselect -> linkdis:chipselect
	wire  [31:0] mm_interconnect_0_linkdis_s1_readdata;     // linkdis:readdata -> mm_interconnect_0:linkdis_s1_readdata
	wire   [1:0] mm_interconnect_0_linkdis_s1_address;      // mm_interconnect_0:linkdis_s1_address -> linkdis:address
	wire         mm_interconnect_0_linkdis_s1_write;        // mm_interconnect_0:linkdis_s1_write -> linkdis:write_n
	wire  [31:0] mm_interconnect_0_linkdis_s1_writedata;    // mm_interconnect_0:linkdis_s1_writedata -> linkdis:writedata
	wire         mm_interconnect_0_linkstart_s1_chipselect; // mm_interconnect_0:linkstart_s1_chipselect -> linkstart:chipselect
	wire  [31:0] mm_interconnect_0_linkstart_s1_readdata;   // linkstart:readdata -> mm_interconnect_0:linkstart_s1_readdata
	wire   [1:0] mm_interconnect_0_linkstart_s1_address;    // mm_interconnect_0:linkstart_s1_address -> linkstart:address
	wire         mm_interconnect_0_linkstart_s1_write;      // mm_interconnect_0:linkstart_s1_write -> linkstart:write_n
	wire  [31:0] mm_interconnect_0_linkstart_s1_writedata;  // mm_interconnect_0:linkstart_s1_writedata -> linkstart:writedata
	wire  [31:0] mm_interconnect_0_rxdata_s1_readdata;      // rxdata:readdata -> mm_interconnect_0:rxdata_s1_readdata
	wire   [1:0] mm_interconnect_0_rxdata_s1_address;       // mm_interconnect_0:rxdata_s1_address -> rxdata:address
	wire  [31:0] mm_interconnect_0_rxflag_s1_readdata;      // rxflag:readdata -> mm_interconnect_0:rxflag_s1_readdata
	wire   [1:0] mm_interconnect_0_rxflag_s1_address;       // mm_interconnect_0:rxflag_s1_address -> rxflag:address
	wire         mm_interconnect_0_txdata_s1_chipselect;    // mm_interconnect_0:txdata_s1_chipselect -> txdata:chipselect
	wire  [31:0] mm_interconnect_0_txdata_s1_readdata;      // txdata:readdata -> mm_interconnect_0:txdata_s1_readdata
	wire   [1:0] mm_interconnect_0_txdata_s1_address;       // mm_interconnect_0:txdata_s1_address -> txdata:address
	wire         mm_interconnect_0_txdata_s1_write;         // mm_interconnect_0:txdata_s1_write -> txdata:write_n
	wire  [31:0] mm_interconnect_0_txdata_s1_writedata;     // mm_interconnect_0:txdata_s1_writedata -> txdata:writedata
	wire         mm_interconnect_0_txflag_s1_chipselect;    // mm_interconnect_0:txflag_s1_chipselect -> txflag:chipselect
	wire  [31:0] mm_interconnect_0_txflag_s1_readdata;      // txflag:readdata -> mm_interconnect_0:txflag_s1_readdata
	wire   [1:0] mm_interconnect_0_txflag_s1_address;       // mm_interconnect_0:txflag_s1_address -> txflag:address
	wire         mm_interconnect_0_txflag_s1_write;         // mm_interconnect_0:txflag_s1_write -> txflag:write_n
	wire  [31:0] mm_interconnect_0_txflag_s1_writedata;     // mm_interconnect_0:txflag_s1_writedata -> txflag:writedata
	wire         mm_interconnect_0_txwrite_s1_chipselect;   // mm_interconnect_0:txwrite_s1_chipselect -> txwrite:chipselect
	wire  [31:0] mm_interconnect_0_txwrite_s1_readdata;     // txwrite:readdata -> mm_interconnect_0:txwrite_s1_readdata
	wire   [1:0] mm_interconnect_0_txwrite_s1_address;      // mm_interconnect_0:txwrite_s1_address -> txwrite:address
	wire         mm_interconnect_0_txwrite_s1_write;        // mm_interconnect_0:txwrite_s1_write -> txwrite:write_n
	wire  [31:0] mm_interconnect_0_txwrite_s1_writedata;    // mm_interconnect_0:txwrite_s1_writedata -> txwrite:writedata
	wire  [31:0] mm_interconnect_0_txrdy_s1_readdata;       // txrdy:readdata -> mm_interconnect_0:txrdy_s1_readdata
	wire   [1:0] mm_interconnect_0_txrdy_s1_address;        // mm_interconnect_0:txrdy_s1_address -> txrdy:address
	wire         mm_interconnect_0_tick_in_s1_chipselect;   // mm_interconnect_0:tick_in_s1_chipselect -> tick_in:chipselect
	wire  [31:0] mm_interconnect_0_tick_in_s1_readdata;     // tick_in:readdata -> mm_interconnect_0:tick_in_s1_readdata
	wire   [1:0] mm_interconnect_0_tick_in_s1_address;      // mm_interconnect_0:tick_in_s1_address -> tick_in:address
	wire         mm_interconnect_0_tick_in_s1_write;        // mm_interconnect_0:tick_in_s1_write -> tick_in:write_n
	wire  [31:0] mm_interconnect_0_tick_in_s1_writedata;    // mm_interconnect_0:tick_in_s1_writedata -> tick_in:writedata
	wire         mm_interconnect_0_time_in_s1_chipselect;   // mm_interconnect_0:time_in_s1_chipselect -> time_in:chipselect
	wire  [31:0] mm_interconnect_0_time_in_s1_readdata;     // time_in:readdata -> mm_interconnect_0:time_in_s1_readdata
	wire   [1:0] mm_interconnect_0_time_in_s1_address;      // mm_interconnect_0:time_in_s1_address -> time_in:address
	wire         mm_interconnect_0_time_in_s1_write;        // mm_interconnect_0:time_in_s1_write -> time_in:write_n
	wire  [31:0] mm_interconnect_0_time_in_s1_writedata;    // mm_interconnect_0:time_in_s1_writedata -> time_in:writedata
	wire  [31:0] mm_interconnect_0_tick_out_s1_readdata;    // tick_out:readdata -> mm_interconnect_0:tick_out_s1_readdata
	wire   [1:0] mm_interconnect_0_tick_out_s1_address;     // mm_interconnect_0:tick_out_s1_address -> tick_out:address
	wire  [31:0] mm_interconnect_0_time_out_s1_readdata;    // time_out:readdata -> mm_interconnect_0:time_out_s1_readdata
	wire   [1:0] mm_interconnect_0_time_out_s1_address;     // mm_interconnect_0:time_out_s1_address -> time_out:address
	wire  [31:0] mm_interconnect_0_txhalff_s1_readdata;     // txhalff:readdata -> mm_interconnect_0:txhalff_s1_readdata
	wire   [1:0] mm_interconnect_0_txhalff_s1_address;      // mm_interconnect_0:txhalff_s1_address -> txhalff:address
	wire  [31:0] mm_interconnect_0_rxhalff_s1_readdata;     // rxhalff:readdata -> mm_interconnect_0:rxhalff_s1_readdata
	wire   [1:0] mm_interconnect_0_rxhalff_s1_address;      // mm_interconnect_0:rxhalff_s1_address -> rxhalff:address
	wire         mm_interconnect_0_rxread_s1_chipselect;    // mm_interconnect_0:rxread_s1_chipselect -> rxread:chipselect
	wire  [31:0] mm_interconnect_0_rxread_s1_readdata;      // rxread:readdata -> mm_interconnect_0:rxread_s1_readdata
	wire   [1:0] mm_interconnect_0_rxread_s1_address;       // mm_interconnect_0:rxread_s1_address -> rxread:address
	wire         mm_interconnect_0_rxread_s1_write;         // mm_interconnect_0:rxread_s1_write -> rxread:write_n
	wire  [31:0] mm_interconnect_0_rxread_s1_writedata;     // mm_interconnect_0:rxread_s1_writedata -> rxread:writedata
	wire  [31:0] mm_interconnect_0_rxvalid_s1_readdata;     // rxvalid:readdata -> mm_interconnect_0:rxvalid_s1_readdata
	wire   [1:0] mm_interconnect_0_rxvalid_s1_address;      // mm_interconnect_0:rxvalid_s1_address -> rxvalid:address
	wire  [31:0] mm_interconnect_0_connecting_s1_readdata;  // connecting:readdata -> mm_interconnect_0:connecting_s1_readdata
	wire   [1:0] mm_interconnect_0_connecting_s1_address;   // mm_interconnect_0:connecting_s1_address -> connecting:address
	wire         mm_interconnect_0_ctrl_in_s1_chipselect;   // mm_interconnect_0:ctrl_in_s1_chipselect -> ctrl_in:chipselect
	wire  [31:0] mm_interconnect_0_ctrl_in_s1_readdata;     // ctrl_in:readdata -> mm_interconnect_0:ctrl_in_s1_readdata
	wire   [1:0] mm_interconnect_0_ctrl_in_s1_address;      // mm_interconnect_0:ctrl_in_s1_address -> ctrl_in:address
	wire         mm_interconnect_0_ctrl_in_s1_write;        // mm_interconnect_0:ctrl_in_s1_write -> ctrl_in:write_n
	wire  [31:0] mm_interconnect_0_ctrl_in_s1_writedata;    // mm_interconnect_0:ctrl_in_s1_writedata -> ctrl_in:writedata
	wire  [31:0] mm_interconnect_0_ctrl_out_s1_readdata;    // ctrl_out:readdata -> mm_interconnect_0:ctrl_out_s1_readdata
	wire   [1:0] mm_interconnect_0_ctrl_out_s1_address;     // mm_interconnect_0:ctrl_out_s1_address -> ctrl_out:address
	wire  [31:0] mm_interconnect_0_errcred_s1_readdata;     // errcred:readdata -> mm_interconnect_0:errcred_s1_readdata
	wire   [1:0] mm_interconnect_0_errcred_s1_address;      // mm_interconnect_0:errcred_s1_address -> errcred:address
	wire  [31:0] mm_interconnect_0_errdisc_s1_readdata;     // errdisc:readdata -> mm_interconnect_0:errdisc_s1_readdata
	wire   [1:0] mm_interconnect_0_errdisc_s1_address;      // mm_interconnect_0:errdisc_s1_address -> errdisc:address
	wire  [31:0] mm_interconnect_0_erresc_s1_readdata;      // erresc:readdata -> mm_interconnect_0:erresc_s1_readdata
	wire   [1:0] mm_interconnect_0_erresc_s1_address;       // mm_interconnect_0:erresc_s1_address -> erresc:address
	wire  [31:0] mm_interconnect_0_errpar_s1_readdata;      // errpar:readdata -> mm_interconnect_0:errpar_s1_readdata
	wire   [1:0] mm_interconnect_0_errpar_s1_address;       // mm_interconnect_0:errpar_s1_address -> errpar:address
	wire  [31:0] mm_interconnect_0_running_s1_readdata;     // running:readdata -> mm_interconnect_0:running_s1_readdata
	wire   [1:0] mm_interconnect_0_running_s1_address;      // mm_interconnect_0:running_s1_address -> running:address
	wire  [31:0] mm_interconnect_0_started_s1_readdata;     // started:readdata -> mm_interconnect_0:started_s1_readdata
	wire   [1:0] mm_interconnect_0_started_s1_address;      // mm_interconnect_0:started_s1_address -> started:address
	wire         mm_interconnect_0_txdivcnt_s1_chipselect;  // mm_interconnect_0:txdivcnt_s1_chipselect -> txdivcnt:chipselect
	wire  [31:0] mm_interconnect_0_txdivcnt_s1_readdata;    // txdivcnt:readdata -> mm_interconnect_0:txdivcnt_s1_readdata
	wire   [1:0] mm_interconnect_0_txdivcnt_s1_address;     // mm_interconnect_0:txdivcnt_s1_address -> txdivcnt:address
	wire         mm_interconnect_0_txdivcnt_s1_write;       // mm_interconnect_0:txdivcnt_s1_write -> txdivcnt:write_n
	wire  [31:0] mm_interconnect_0_txdivcnt_s1_writedata;   // mm_interconnect_0:txdivcnt_s1_writedata -> txdivcnt:writedata
	wire         rst_controller_reset_out_reset;            // rst_controller:reset_out -> [autostart:reset_n, connecting:reset_n, ctrl_in:reset_n, ctrl_out:reset_n, errcred:reset_n, errdisc:reset_n, erresc:reset_n, errpar:reset_n, linkdis:reset_n, linkstart:reset_n, mm_interconnect_0:autostart_reset_reset_bridge_in_reset_reset, running:reset_n, rxdata:reset_n, rxflag:reset_n, rxhalff:reset_n, rxread:reset_n, rxvalid:reset_n, started:reset_n, tick_in:reset_n, tick_out:reset_n, time_in:reset_n, time_out:reset_n, txdata:reset_n, txdivcnt:reset_n, txflag:reset_n, txhalff:reset_n, txrdy:reset_n, txwrite:reset_n]
	wire         rst_controller_001_reset_out_reset;        // rst_controller_001:reset_out -> mm_interconnect_0:hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset
	wire         hps_0_h2f_reset_reset;                     // hps_0:h2f_rst_n -> rst_controller_001:reset_in0

	spw_light_autostart autostart (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_autostart_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_autostart_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_autostart_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_autostart_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_autostart_s1_readdata),   //                    .readdata
		.out_port   (autostart_external_connection_export)       // external_connection.export
	);

	spw_light_connecting connecting (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_connecting_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_connecting_s1_readdata), //                    .readdata
		.in_port  (connecting_external_connection_export)     // external_connection.export
	);

	spw_light_ctrl_in ctrl_in (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_ctrl_in_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ctrl_in_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ctrl_in_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ctrl_in_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ctrl_in_s1_readdata),   //                    .readdata
		.out_port   (ctrl_in_external_connection_export)       // external_connection.export
	);

	spw_light_ctrl_out ctrl_out (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_ctrl_out_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_ctrl_out_s1_readdata), //                    .readdata
		.in_port  (ctrl_out_external_connection_export)     // external_connection.export
	);

	spw_light_connecting errcred (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_errcred_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_errcred_s1_readdata), //                    .readdata
		.in_port  (errcred_external_connection_export)     // external_connection.export
	);

	spw_light_connecting errdisc (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_errdisc_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_errdisc_s1_readdata), //                    .readdata
		.in_port  (errdisc_external_connection_export)     // external_connection.export
	);

	spw_light_connecting erresc (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_erresc_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_erresc_s1_readdata), //                    .readdata
		.in_port  (erresc_external_connection_export)     // external_connection.export
	);

	spw_light_connecting errpar (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_errpar_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_errpar_s1_readdata), //                    .readdata
		.in_port  (errpar_external_connection_export)     // external_connection.export
	);

	spw_light_hps_0 #(
		.F2S_Width (0),
		.S2F_Width (1)
	) hps_0 (
		.mem_a       (memory_mem_a),                 //         memory.mem_a
		.mem_ba      (memory_mem_ba),                //               .mem_ba
		.mem_ck      (memory_mem_ck),                //               .mem_ck
		.mem_ck_n    (memory_mem_ck_n),              //               .mem_ck_n
		.mem_cke     (memory_mem_cke),               //               .mem_cke
		.mem_cs_n    (memory_mem_cs_n),              //               .mem_cs_n
		.mem_ras_n   (memory_mem_ras_n),             //               .mem_ras_n
		.mem_cas_n   (memory_mem_cas_n),             //               .mem_cas_n
		.mem_we_n    (memory_mem_we_n),              //               .mem_we_n
		.mem_reset_n (memory_mem_reset_n),           //               .mem_reset_n
		.mem_dq      (memory_mem_dq),                //               .mem_dq
		.mem_dqs     (memory_mem_dqs),               //               .mem_dqs
		.mem_dqs_n   (memory_mem_dqs_n),             //               .mem_dqs_n
		.mem_odt     (memory_mem_odt),               //               .mem_odt
		.mem_dm      (memory_mem_dm),                //               .mem_dm
		.oct_rzqin   (memory_oct_rzqin),             //               .oct_rzqin
		.h2f_rst_n   (hps_0_h2f_reset_reset),        //      h2f_reset.reset_n
		.h2f_axi_clk (clk_clk),                      //  h2f_axi_clock.clk
		.h2f_AWID    (hps_0_h2f_axi_master_awid),    // h2f_axi_master.awid
		.h2f_AWADDR  (hps_0_h2f_axi_master_awaddr),  //               .awaddr
		.h2f_AWLEN   (hps_0_h2f_axi_master_awlen),   //               .awlen
		.h2f_AWSIZE  (hps_0_h2f_axi_master_awsize),  //               .awsize
		.h2f_AWBURST (hps_0_h2f_axi_master_awburst), //               .awburst
		.h2f_AWLOCK  (hps_0_h2f_axi_master_awlock),  //               .awlock
		.h2f_AWCACHE (hps_0_h2f_axi_master_awcache), //               .awcache
		.h2f_AWPROT  (hps_0_h2f_axi_master_awprot),  //               .awprot
		.h2f_AWVALID (hps_0_h2f_axi_master_awvalid), //               .awvalid
		.h2f_AWREADY (hps_0_h2f_axi_master_awready), //               .awready
		.h2f_WID     (hps_0_h2f_axi_master_wid),     //               .wid
		.h2f_WDATA   (hps_0_h2f_axi_master_wdata),   //               .wdata
		.h2f_WSTRB   (hps_0_h2f_axi_master_wstrb),   //               .wstrb
		.h2f_WLAST   (hps_0_h2f_axi_master_wlast),   //               .wlast
		.h2f_WVALID  (hps_0_h2f_axi_master_wvalid),  //               .wvalid
		.h2f_WREADY  (hps_0_h2f_axi_master_wready),  //               .wready
		.h2f_BID     (hps_0_h2f_axi_master_bid),     //               .bid
		.h2f_BRESP   (hps_0_h2f_axi_master_bresp),   //               .bresp
		.h2f_BVALID  (hps_0_h2f_axi_master_bvalid),  //               .bvalid
		.h2f_BREADY  (hps_0_h2f_axi_master_bready),  //               .bready
		.h2f_ARID    (hps_0_h2f_axi_master_arid),    //               .arid
		.h2f_ARADDR  (hps_0_h2f_axi_master_araddr),  //               .araddr
		.h2f_ARLEN   (hps_0_h2f_axi_master_arlen),   //               .arlen
		.h2f_ARSIZE  (hps_0_h2f_axi_master_arsize),  //               .arsize
		.h2f_ARBURST (hps_0_h2f_axi_master_arburst), //               .arburst
		.h2f_ARLOCK  (hps_0_h2f_axi_master_arlock),  //               .arlock
		.h2f_ARCACHE (hps_0_h2f_axi_master_arcache), //               .arcache
		.h2f_ARPROT  (hps_0_h2f_axi_master_arprot),  //               .arprot
		.h2f_ARVALID (hps_0_h2f_axi_master_arvalid), //               .arvalid
		.h2f_ARREADY (hps_0_h2f_axi_master_arready), //               .arready
		.h2f_RID     (hps_0_h2f_axi_master_rid),     //               .rid
		.h2f_RDATA   (hps_0_h2f_axi_master_rdata),   //               .rdata
		.h2f_RRESP   (hps_0_h2f_axi_master_rresp),   //               .rresp
		.h2f_RLAST   (hps_0_h2f_axi_master_rlast),   //               .rlast
		.h2f_RVALID  (hps_0_h2f_axi_master_rvalid),  //               .rvalid
		.h2f_RREADY  (hps_0_h2f_axi_master_rready)   //               .rready
	);

	spw_light_autostart linkdis (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_linkdis_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_linkdis_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_linkdis_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_linkdis_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_linkdis_s1_readdata),   //                    .readdata
		.out_port   (linkdis_external_connection_export)       // external_connection.export
	);

	spw_light_autostart linkstart (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_linkstart_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_linkstart_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_linkstart_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_linkstart_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_linkstart_s1_readdata),   //                    .readdata
		.out_port   (linkstart_external_connection_export)       // external_connection.export
	);

	spw_light_pll_0 pll_0 (
		.refclk   (clk_clk),             //  refclk.clk
		.rst      (~reset_reset_n),      //   reset.reset
		.outclk_0 (pll_0_outclk0_clk),   // outclk0.clk
		.locked   (pll_0_locked_export)  //  locked.export
	);

	spw_light_connecting running (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_running_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_running_s1_readdata), //                    .readdata
		.in_port  (running_external_connection_export)     // external_connection.export
	);

	spw_light_rxdata rxdata (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_rxdata_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_rxdata_s1_readdata), //                    .readdata
		.in_port  (rxdata_external_connection_export)     // external_connection.export
	);

	spw_light_connecting rxflag (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_rxflag_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_rxflag_s1_readdata), //                    .readdata
		.in_port  (rxflag_external_connection_export)     // external_connection.export
	);

	spw_light_connecting rxhalff (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_rxhalff_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_rxhalff_s1_readdata), //                    .readdata
		.in_port  (rxhalff_external_connection_export)     // external_connection.export
	);

	spw_light_autostart rxread (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_rxread_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_rxread_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_rxread_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_rxread_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_rxread_s1_readdata),   //                    .readdata
		.out_port   (rxread_external_connection_export)       // external_connection.export
	);

	spw_light_connecting rxvalid (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_rxvalid_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_rxvalid_s1_readdata), //                    .readdata
		.in_port  (rxvalid_external_connection_export)     // external_connection.export
	);

	spw_light_connecting started (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_started_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_started_s1_readdata), //                    .readdata
		.in_port  (started_external_connection_export)     // external_connection.export
	);

	spw_light_autostart tick_in (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_tick_in_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_tick_in_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_tick_in_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_tick_in_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_tick_in_s1_readdata),   //                    .readdata
		.out_port   (tick_in_external_connection_export)       // external_connection.export
	);

	spw_light_connecting tick_out (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_tick_out_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_tick_out_s1_readdata), //                    .readdata
		.in_port  (tick_out_external_connection_export)     // external_connection.export
	);

	spw_light_time_in time_in (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_time_in_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_time_in_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_time_in_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_time_in_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_time_in_s1_readdata),   //                    .readdata
		.out_port   (time_in_external_connection_export)       // external_connection.export
	);

	spw_light_time_out time_out (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_time_out_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_time_out_s1_readdata), //                    .readdata
		.in_port  (time_out_external_connection_export)     // external_connection.export
	);

	spw_light_txdata txdata (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_txdata_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_txdata_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_txdata_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_txdata_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_txdata_s1_readdata),   //                    .readdata
		.out_port   (txdata_external_connection_export)       // external_connection.export
	);

	spw_light_txdata txdivcnt (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_txdivcnt_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_txdivcnt_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_txdivcnt_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_txdivcnt_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_txdivcnt_s1_readdata),   //                    .readdata
		.out_port   (txdivcnt_external_connection_export)       // external_connection.export
	);

	spw_light_autostart txflag (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_txflag_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_txflag_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_txflag_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_txflag_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_txflag_s1_readdata),   //                    .readdata
		.out_port   (txflag_external_connection_export)       // external_connection.export
	);

	spw_light_connecting txhalff (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_txhalff_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_txhalff_s1_readdata), //                    .readdata
		.in_port  (txhalff_external_connection_export)     // external_connection.export
	);

	spw_light_connecting txrdy (
		.clk      (clk_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_txrdy_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_txrdy_s1_readdata), //                    .readdata
		.in_port  (txrdy_external_connection_export)     // external_connection.export
	);

	spw_light_autostart txwrite (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_txwrite_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_txwrite_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_txwrite_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_txwrite_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_txwrite_s1_readdata),   //                    .readdata
		.out_port   (txwrite_external_connection_export)       // external_connection.export
	);

	spw_light_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_h2f_axi_master_awid                                        (hps_0_h2f_axi_master_awid),                 //                                       hps_0_h2f_axi_master.awid
		.hps_0_h2f_axi_master_awaddr                                      (hps_0_h2f_axi_master_awaddr),               //                                                           .awaddr
		.hps_0_h2f_axi_master_awlen                                       (hps_0_h2f_axi_master_awlen),                //                                                           .awlen
		.hps_0_h2f_axi_master_awsize                                      (hps_0_h2f_axi_master_awsize),               //                                                           .awsize
		.hps_0_h2f_axi_master_awburst                                     (hps_0_h2f_axi_master_awburst),              //                                                           .awburst
		.hps_0_h2f_axi_master_awlock                                      (hps_0_h2f_axi_master_awlock),               //                                                           .awlock
		.hps_0_h2f_axi_master_awcache                                     (hps_0_h2f_axi_master_awcache),              //                                                           .awcache
		.hps_0_h2f_axi_master_awprot                                      (hps_0_h2f_axi_master_awprot),               //                                                           .awprot
		.hps_0_h2f_axi_master_awvalid                                     (hps_0_h2f_axi_master_awvalid),              //                                                           .awvalid
		.hps_0_h2f_axi_master_awready                                     (hps_0_h2f_axi_master_awready),              //                                                           .awready
		.hps_0_h2f_axi_master_wid                                         (hps_0_h2f_axi_master_wid),                  //                                                           .wid
		.hps_0_h2f_axi_master_wdata                                       (hps_0_h2f_axi_master_wdata),                //                                                           .wdata
		.hps_0_h2f_axi_master_wstrb                                       (hps_0_h2f_axi_master_wstrb),                //                                                           .wstrb
		.hps_0_h2f_axi_master_wlast                                       (hps_0_h2f_axi_master_wlast),                //                                                           .wlast
		.hps_0_h2f_axi_master_wvalid                                      (hps_0_h2f_axi_master_wvalid),               //                                                           .wvalid
		.hps_0_h2f_axi_master_wready                                      (hps_0_h2f_axi_master_wready),               //                                                           .wready
		.hps_0_h2f_axi_master_bid                                         (hps_0_h2f_axi_master_bid),                  //                                                           .bid
		.hps_0_h2f_axi_master_bresp                                       (hps_0_h2f_axi_master_bresp),                //                                                           .bresp
		.hps_0_h2f_axi_master_bvalid                                      (hps_0_h2f_axi_master_bvalid),               //                                                           .bvalid
		.hps_0_h2f_axi_master_bready                                      (hps_0_h2f_axi_master_bready),               //                                                           .bready
		.hps_0_h2f_axi_master_arid                                        (hps_0_h2f_axi_master_arid),                 //                                                           .arid
		.hps_0_h2f_axi_master_araddr                                      (hps_0_h2f_axi_master_araddr),               //                                                           .araddr
		.hps_0_h2f_axi_master_arlen                                       (hps_0_h2f_axi_master_arlen),                //                                                           .arlen
		.hps_0_h2f_axi_master_arsize                                      (hps_0_h2f_axi_master_arsize),               //                                                           .arsize
		.hps_0_h2f_axi_master_arburst                                     (hps_0_h2f_axi_master_arburst),              //                                                           .arburst
		.hps_0_h2f_axi_master_arlock                                      (hps_0_h2f_axi_master_arlock),               //                                                           .arlock
		.hps_0_h2f_axi_master_arcache                                     (hps_0_h2f_axi_master_arcache),              //                                                           .arcache
		.hps_0_h2f_axi_master_arprot                                      (hps_0_h2f_axi_master_arprot),               //                                                           .arprot
		.hps_0_h2f_axi_master_arvalid                                     (hps_0_h2f_axi_master_arvalid),              //                                                           .arvalid
		.hps_0_h2f_axi_master_arready                                     (hps_0_h2f_axi_master_arready),              //                                                           .arready
		.hps_0_h2f_axi_master_rid                                         (hps_0_h2f_axi_master_rid),                  //                                                           .rid
		.hps_0_h2f_axi_master_rdata                                       (hps_0_h2f_axi_master_rdata),                //                                                           .rdata
		.hps_0_h2f_axi_master_rresp                                       (hps_0_h2f_axi_master_rresp),                //                                                           .rresp
		.hps_0_h2f_axi_master_rlast                                       (hps_0_h2f_axi_master_rlast),                //                                                           .rlast
		.hps_0_h2f_axi_master_rvalid                                      (hps_0_h2f_axi_master_rvalid),               //                                                           .rvalid
		.hps_0_h2f_axi_master_rready                                      (hps_0_h2f_axi_master_rready),               //                                                           .rready
		.clk_0_clk_clk                                                    (clk_clk),                                   //                                                  clk_0_clk.clk
		.autostart_reset_reset_bridge_in_reset_reset                      (rst_controller_reset_out_reset),            //                      autostart_reset_reset_bridge_in_reset.reset
		.hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),        // hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.autostart_s1_address                                             (mm_interconnect_0_autostart_s1_address),    //                                               autostart_s1.address
		.autostart_s1_write                                               (mm_interconnect_0_autostart_s1_write),      //                                                           .write
		.autostart_s1_readdata                                            (mm_interconnect_0_autostart_s1_readdata),   //                                                           .readdata
		.autostart_s1_writedata                                           (mm_interconnect_0_autostart_s1_writedata),  //                                                           .writedata
		.autostart_s1_chipselect                                          (mm_interconnect_0_autostart_s1_chipselect), //                                                           .chipselect
		.connecting_s1_address                                            (mm_interconnect_0_connecting_s1_address),   //                                              connecting_s1.address
		.connecting_s1_readdata                                           (mm_interconnect_0_connecting_s1_readdata),  //                                                           .readdata
		.ctrl_in_s1_address                                               (mm_interconnect_0_ctrl_in_s1_address),      //                                                 ctrl_in_s1.address
		.ctrl_in_s1_write                                                 (mm_interconnect_0_ctrl_in_s1_write),        //                                                           .write
		.ctrl_in_s1_readdata                                              (mm_interconnect_0_ctrl_in_s1_readdata),     //                                                           .readdata
		.ctrl_in_s1_writedata                                             (mm_interconnect_0_ctrl_in_s1_writedata),    //                                                           .writedata
		.ctrl_in_s1_chipselect                                            (mm_interconnect_0_ctrl_in_s1_chipselect),   //                                                           .chipselect
		.ctrl_out_s1_address                                              (mm_interconnect_0_ctrl_out_s1_address),     //                                                ctrl_out_s1.address
		.ctrl_out_s1_readdata                                             (mm_interconnect_0_ctrl_out_s1_readdata),    //                                                           .readdata
		.errcred_s1_address                                               (mm_interconnect_0_errcred_s1_address),      //                                                 errcred_s1.address
		.errcred_s1_readdata                                              (mm_interconnect_0_errcred_s1_readdata),     //                                                           .readdata
		.errdisc_s1_address                                               (mm_interconnect_0_errdisc_s1_address),      //                                                 errdisc_s1.address
		.errdisc_s1_readdata                                              (mm_interconnect_0_errdisc_s1_readdata),     //                                                           .readdata
		.erresc_s1_address                                                (mm_interconnect_0_erresc_s1_address),       //                                                  erresc_s1.address
		.erresc_s1_readdata                                               (mm_interconnect_0_erresc_s1_readdata),      //                                                           .readdata
		.errpar_s1_address                                                (mm_interconnect_0_errpar_s1_address),       //                                                  errpar_s1.address
		.errpar_s1_readdata                                               (mm_interconnect_0_errpar_s1_readdata),      //                                                           .readdata
		.linkdis_s1_address                                               (mm_interconnect_0_linkdis_s1_address),      //                                                 linkdis_s1.address
		.linkdis_s1_write                                                 (mm_interconnect_0_linkdis_s1_write),        //                                                           .write
		.linkdis_s1_readdata                                              (mm_interconnect_0_linkdis_s1_readdata),     //                                                           .readdata
		.linkdis_s1_writedata                                             (mm_interconnect_0_linkdis_s1_writedata),    //                                                           .writedata
		.linkdis_s1_chipselect                                            (mm_interconnect_0_linkdis_s1_chipselect),   //                                                           .chipselect
		.linkstart_s1_address                                             (mm_interconnect_0_linkstart_s1_address),    //                                               linkstart_s1.address
		.linkstart_s1_write                                               (mm_interconnect_0_linkstart_s1_write),      //                                                           .write
		.linkstart_s1_readdata                                            (mm_interconnect_0_linkstart_s1_readdata),   //                                                           .readdata
		.linkstart_s1_writedata                                           (mm_interconnect_0_linkstart_s1_writedata),  //                                                           .writedata
		.linkstart_s1_chipselect                                          (mm_interconnect_0_linkstart_s1_chipselect), //                                                           .chipselect
		.running_s1_address                                               (mm_interconnect_0_running_s1_address),      //                                                 running_s1.address
		.running_s1_readdata                                              (mm_interconnect_0_running_s1_readdata),     //                                                           .readdata
		.rxdata_s1_address                                                (mm_interconnect_0_rxdata_s1_address),       //                                                  rxdata_s1.address
		.rxdata_s1_readdata                                               (mm_interconnect_0_rxdata_s1_readdata),      //                                                           .readdata
		.rxflag_s1_address                                                (mm_interconnect_0_rxflag_s1_address),       //                                                  rxflag_s1.address
		.rxflag_s1_readdata                                               (mm_interconnect_0_rxflag_s1_readdata),      //                                                           .readdata
		.rxhalff_s1_address                                               (mm_interconnect_0_rxhalff_s1_address),      //                                                 rxhalff_s1.address
		.rxhalff_s1_readdata                                              (mm_interconnect_0_rxhalff_s1_readdata),     //                                                           .readdata
		.rxread_s1_address                                                (mm_interconnect_0_rxread_s1_address),       //                                                  rxread_s1.address
		.rxread_s1_write                                                  (mm_interconnect_0_rxread_s1_write),         //                                                           .write
		.rxread_s1_readdata                                               (mm_interconnect_0_rxread_s1_readdata),      //                                                           .readdata
		.rxread_s1_writedata                                              (mm_interconnect_0_rxread_s1_writedata),     //                                                           .writedata
		.rxread_s1_chipselect                                             (mm_interconnect_0_rxread_s1_chipselect),    //                                                           .chipselect
		.rxvalid_s1_address                                               (mm_interconnect_0_rxvalid_s1_address),      //                                                 rxvalid_s1.address
		.rxvalid_s1_readdata                                              (mm_interconnect_0_rxvalid_s1_readdata),     //                                                           .readdata
		.started_s1_address                                               (mm_interconnect_0_started_s1_address),      //                                                 started_s1.address
		.started_s1_readdata                                              (mm_interconnect_0_started_s1_readdata),     //                                                           .readdata
		.tick_in_s1_address                                               (mm_interconnect_0_tick_in_s1_address),      //                                                 tick_in_s1.address
		.tick_in_s1_write                                                 (mm_interconnect_0_tick_in_s1_write),        //                                                           .write
		.tick_in_s1_readdata                                              (mm_interconnect_0_tick_in_s1_readdata),     //                                                           .readdata
		.tick_in_s1_writedata                                             (mm_interconnect_0_tick_in_s1_writedata),    //                                                           .writedata
		.tick_in_s1_chipselect                                            (mm_interconnect_0_tick_in_s1_chipselect),   //                                                           .chipselect
		.tick_out_s1_address                                              (mm_interconnect_0_tick_out_s1_address),     //                                                tick_out_s1.address
		.tick_out_s1_readdata                                             (mm_interconnect_0_tick_out_s1_readdata),    //                                                           .readdata
		.time_in_s1_address                                               (mm_interconnect_0_time_in_s1_address),      //                                                 time_in_s1.address
		.time_in_s1_write                                                 (mm_interconnect_0_time_in_s1_write),        //                                                           .write
		.time_in_s1_readdata                                              (mm_interconnect_0_time_in_s1_readdata),     //                                                           .readdata
		.time_in_s1_writedata                                             (mm_interconnect_0_time_in_s1_writedata),    //                                                           .writedata
		.time_in_s1_chipselect                                            (mm_interconnect_0_time_in_s1_chipselect),   //                                                           .chipselect
		.time_out_s1_address                                              (mm_interconnect_0_time_out_s1_address),     //                                                time_out_s1.address
		.time_out_s1_readdata                                             (mm_interconnect_0_time_out_s1_readdata),    //                                                           .readdata
		.txdata_s1_address                                                (mm_interconnect_0_txdata_s1_address),       //                                                  txdata_s1.address
		.txdata_s1_write                                                  (mm_interconnect_0_txdata_s1_write),         //                                                           .write
		.txdata_s1_readdata                                               (mm_interconnect_0_txdata_s1_readdata),      //                                                           .readdata
		.txdata_s1_writedata                                              (mm_interconnect_0_txdata_s1_writedata),     //                                                           .writedata
		.txdata_s1_chipselect                                             (mm_interconnect_0_txdata_s1_chipselect),    //                                                           .chipselect
		.txdivcnt_s1_address                                              (mm_interconnect_0_txdivcnt_s1_address),     //                                                txdivcnt_s1.address
		.txdivcnt_s1_write                                                (mm_interconnect_0_txdivcnt_s1_write),       //                                                           .write
		.txdivcnt_s1_readdata                                             (mm_interconnect_0_txdivcnt_s1_readdata),    //                                                           .readdata
		.txdivcnt_s1_writedata                                            (mm_interconnect_0_txdivcnt_s1_writedata),   //                                                           .writedata
		.txdivcnt_s1_chipselect                                           (mm_interconnect_0_txdivcnt_s1_chipselect),  //                                                           .chipselect
		.txflag_s1_address                                                (mm_interconnect_0_txflag_s1_address),       //                                                  txflag_s1.address
		.txflag_s1_write                                                  (mm_interconnect_0_txflag_s1_write),         //                                                           .write
		.txflag_s1_readdata                                               (mm_interconnect_0_txflag_s1_readdata),      //                                                           .readdata
		.txflag_s1_writedata                                              (mm_interconnect_0_txflag_s1_writedata),     //                                                           .writedata
		.txflag_s1_chipselect                                             (mm_interconnect_0_txflag_s1_chipselect),    //                                                           .chipselect
		.txhalff_s1_address                                               (mm_interconnect_0_txhalff_s1_address),      //                                                 txhalff_s1.address
		.txhalff_s1_readdata                                              (mm_interconnect_0_txhalff_s1_readdata),     //                                                           .readdata
		.txrdy_s1_address                                                 (mm_interconnect_0_txrdy_s1_address),        //                                                   txrdy_s1.address
		.txrdy_s1_readdata                                                (mm_interconnect_0_txrdy_s1_readdata),       //                                                           .readdata
		.txwrite_s1_address                                               (mm_interconnect_0_txwrite_s1_address),      //                                                 txwrite_s1.address
		.txwrite_s1_write                                                 (mm_interconnect_0_txwrite_s1_write),        //                                                           .write
		.txwrite_s1_readdata                                              (mm_interconnect_0_txwrite_s1_readdata),     //                                                           .readdata
		.txwrite_s1_writedata                                             (mm_interconnect_0_txwrite_s1_writedata),    //                                                           .writedata
		.txwrite_s1_chipselect                                            (mm_interconnect_0_txwrite_s1_chipselect)    //                                                           .chipselect
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~hps_0_h2f_reset_reset),             // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
