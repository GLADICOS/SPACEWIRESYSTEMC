-- jaxa.vhd

-- Generated using ACDS version 17.1 593

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity jaxa is
	port (
		autostart_external_connection_export                   : out   std_logic;                                        --                   autostart_external_connection.export
		clk_clk                                                : in    std_logic                     := '0';             --                                             clk.clk
		controlflagsin_external_connection_export              : out   std_logic_vector(1 downto 0);                     --              controlflagsin_external_connection.export
		controlflagsout_external_connection_export             : in    std_logic_vector(1 downto 0)  := (others => '0'); --             controlflagsout_external_connection.export
		creditcount_external_connection_export                 : in    std_logic_vector(5 downto 0)  := (others => '0'); --                 creditcount_external_connection.export
		errorstatus_external_connection_export                 : in    std_logic_vector(7 downto 0)  := (others => '0'); --                 errorstatus_external_connection.export
		linkdisable_external_connection_export                 : out   std_logic;                                        --                 linkdisable_external_connection.export
		linkstart_external_connection_export                   : out   std_logic;                                        --                   linkstart_external_connection.export
		linkstatus_external_connection_export                  : in    std_logic_vector(15 downto 0) := (others => '0'); --                  linkstatus_external_connection.export
		memory_mem_a                                           : out   std_logic_vector(12 downto 0);                    --                                          memory.mem_a
		memory_mem_ba                                          : out   std_logic_vector(2 downto 0);                     --                                                .mem_ba
		memory_mem_ck                                          : out   std_logic;                                        --                                                .mem_ck
		memory_mem_ck_n                                        : out   std_logic;                                        --                                                .mem_ck_n
		memory_mem_cke                                         : out   std_logic;                                        --                                                .mem_cke
		memory_mem_cs_n                                        : out   std_logic;                                        --                                                .mem_cs_n
		memory_mem_ras_n                                       : out   std_logic;                                        --                                                .mem_ras_n
		memory_mem_cas_n                                       : out   std_logic;                                        --                                                .mem_cas_n
		memory_mem_we_n                                        : out   std_logic;                                        --                                                .mem_we_n
		memory_mem_reset_n                                     : out   std_logic;                                        --                                                .mem_reset_n
		memory_mem_dq                                          : inout std_logic_vector(7 downto 0)  := (others => '0'); --                                                .mem_dq
		memory_mem_dqs                                         : inout std_logic                     := '0';             --                                                .mem_dqs
		memory_mem_dqs_n                                       : inout std_logic                     := '0';             --                                                .mem_dqs_n
		memory_mem_odt                                         : out   std_logic;                                        --                                                .mem_odt
		memory_mem_dm                                          : out   std_logic;                                        --                                                .mem_dm
		memory_oct_rzqin                                       : in    std_logic                     := '0';             --                                                .oct_rzqin
		outstandingcount_external_connection_export            : in    std_logic_vector(5 downto 0)  := (others => '0'); --            outstandingcount_external_connection.export
		pll_0_outclk0_clk                                      : out   std_logic;                                        --                                   pll_0_outclk0.clk
		receiveactivity_external_connection_export             : in    std_logic                     := '0';             --             receiveactivity_external_connection.export
		receiveclock_external_connection_export                : out   std_logic;                                        --                receiveclock_external_connection.export
		receivefifodatacount_external_connection_export        : in    std_logic                     := '0';             --        receivefifodatacount_external_connection.export
		receivefifodataout_external_connection_export          : in    std_logic_vector(8 downto 0)  := (others => '0'); --          receivefifodataout_external_connection.export
		receivefifoempty_external_connection_export            : in    std_logic                     := '0';             --            receivefifoempty_external_connection.export
		receivefifofull_external_connection_export             : in    std_logic                     := '0';             --             receivefifofull_external_connection.export
		receivefiforeadenable_external_connection_export       : out   std_logic;                                        --       receivefiforeadenable_external_connection.export
		spacewiredatain_external_connection_export             : out   std_logic;                                        --             spacewiredatain_external_connection.export
		spacewiredataout_external_connection_export            : in    std_logic                     := '0';             --            spacewiredataout_external_connection.export
		spacewirestrobein_external_connection_export           : out   std_logic;                                        --           spacewirestrobein_external_connection.export
		spacewirestrobeout_external_connection_export          : in    std_logic                     := '0';             --          spacewirestrobeout_external_connection.export
		statisticalinformation_0_external_connection_export    : in    std_logic_vector(31 downto 0) := (others => '0'); --    statisticalinformation_0_external_connection.export
		statisticalinformation_1_external_connection_export    : in    std_logic_vector(31 downto 0) := (others => '0'); --    statisticalinformation_1_external_connection.export
		statisticalinformation_2_external_connection_export    : in    std_logic_vector(31 downto 0) := (others => '0'); --    statisticalinformation_2_external_connection.export
		statisticalinformation_3_external_connection_export    : in    std_logic_vector(31 downto 0) := (others => '0'); --    statisticalinformation_3_external_connection.export
		statisticalinformation_4_external_connection_export    : in    std_logic_vector(31 downto 0) := (others => '0'); --    statisticalinformation_4_external_connection.export
		statisticalinformation_5_external_connection_export    : in    std_logic_vector(31 downto 0) := (others => '0'); --    statisticalinformation_5_external_connection.export
		statisticalinformation_6_external_connection_export    : in    std_logic_vector(31 downto 0) := (others => '0'); --    statisticalinformation_6_external_connection.export
		statisticalinformation_7_external_connection_export    : in    std_logic_vector(31 downto 0) := (others => '0'); --    statisticalinformation_7_external_connection.export
		statisticalinformationclear_external_connection_export : out   std_logic;                                        -- statisticalinformationclear_external_connection.export
		tickin_external_connection_export                      : out   std_logic;                                        --                      tickin_external_connection.export
		tickout_external_connection_export                     : in    std_logic                     := '0';             --                     tickout_external_connection.export
		timein_external_connection_export                      : out   std_logic_vector(5 downto 0);                     --                      timein_external_connection.export
		timeout_external_connection_export                     : in    std_logic_vector(5 downto 0)  := (others => '0'); --                     timeout_external_connection.export
		transmitactivity_external_connection_export            : in    std_logic                     := '0';             --            transmitactivity_external_connection.export
		transmitclock_external_connection_export               : out   std_logic;                                        --               transmitclock_external_connection.export
		transmitclockdividevalue_external_connection_export    : out   std_logic_vector(5 downto 0);                     --    transmitclockdividevalue_external_connection.export
		transmitfifodatacount_external_connection_export       : in    std_logic_vector(5 downto 0)  := (others => '0'); --       transmitfifodatacount_external_connection.export
		transmitfifodatain_external_connection_export          : out   std_logic_vector(8 downto 0);                     --          transmitfifodatain_external_connection.export
		transmitfifofull_external_connection_export            : in    std_logic                     := '0';             --            transmitfifofull_external_connection.export
		transmitfifowriteenable_external_connection_export     : out   std_logic                                         --     transmitfifowriteenable_external_connection.export
	);
end entity jaxa;

architecture rtl of jaxa is
	component jaxa_autoStart is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic                                         -- export
		);
	end component jaxa_autoStart;

	component jaxa_controlFlagsIn is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(1 downto 0)                      -- export
		);
	end component jaxa_controlFlagsIn;

	component jaxa_controlFlagsOut is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(1 downto 0)  := (others => 'X')  -- export
		);
	end component jaxa_controlFlagsOut;

	component jaxa_creditCount is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(5 downto 0)  := (others => 'X')  -- export
		);
	end component jaxa_creditCount;

	component jaxa_errorStatus is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- export
		);
	end component jaxa_errorStatus;

	component jaxa_hps_0 is
		generic (
			F2S_Width : integer := 2;
			S2F_Width : integer := 2
		);
		port (
			mem_a       : out   std_logic_vector(12 downto 0);                    -- mem_a
			mem_ba      : out   std_logic_vector(2 downto 0);                     -- mem_ba
			mem_ck      : out   std_logic;                                        -- mem_ck
			mem_ck_n    : out   std_logic;                                        -- mem_ck_n
			mem_cke     : out   std_logic;                                        -- mem_cke
			mem_cs_n    : out   std_logic;                                        -- mem_cs_n
			mem_ras_n   : out   std_logic;                                        -- mem_ras_n
			mem_cas_n   : out   std_logic;                                        -- mem_cas_n
			mem_we_n    : out   std_logic;                                        -- mem_we_n
			mem_reset_n : out   std_logic;                                        -- mem_reset_n
			mem_dq      : inout std_logic_vector(7 downto 0)  := (others => 'X'); -- mem_dq
			mem_dqs     : inout std_logic                     := 'X';             -- mem_dqs
			mem_dqs_n   : inout std_logic                     := 'X';             -- mem_dqs_n
			mem_odt     : out   std_logic;                                        -- mem_odt
			mem_dm      : out   std_logic;                                        -- mem_dm
			oct_rzqin   : in    std_logic                     := 'X';             -- oct_rzqin
			h2f_rst_n   : out   std_logic;                                        -- reset_n
			h2f_axi_clk : in    std_logic                     := 'X';             -- clk
			h2f_AWID    : out   std_logic_vector(11 downto 0);                    -- awid
			h2f_AWADDR  : out   std_logic_vector(29 downto 0);                    -- awaddr
			h2f_AWLEN   : out   std_logic_vector(3 downto 0);                     -- awlen
			h2f_AWSIZE  : out   std_logic_vector(2 downto 0);                     -- awsize
			h2f_AWBURST : out   std_logic_vector(1 downto 0);                     -- awburst
			h2f_AWLOCK  : out   std_logic_vector(1 downto 0);                     -- awlock
			h2f_AWCACHE : out   std_logic_vector(3 downto 0);                     -- awcache
			h2f_AWPROT  : out   std_logic_vector(2 downto 0);                     -- awprot
			h2f_AWVALID : out   std_logic;                                        -- awvalid
			h2f_AWREADY : in    std_logic                     := 'X';             -- awready
			h2f_WID     : out   std_logic_vector(11 downto 0);                    -- wid
			h2f_WDATA   : out   std_logic_vector(31 downto 0);                    -- wdata
			h2f_WSTRB   : out   std_logic_vector(3 downto 0);                     -- wstrb
			h2f_WLAST   : out   std_logic;                                        -- wlast
			h2f_WVALID  : out   std_logic;                                        -- wvalid
			h2f_WREADY  : in    std_logic                     := 'X';             -- wready
			h2f_BID     : in    std_logic_vector(11 downto 0) := (others => 'X'); -- bid
			h2f_BRESP   : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			h2f_BVALID  : in    std_logic                     := 'X';             -- bvalid
			h2f_BREADY  : out   std_logic;                                        -- bready
			h2f_ARID    : out   std_logic_vector(11 downto 0);                    -- arid
			h2f_ARADDR  : out   std_logic_vector(29 downto 0);                    -- araddr
			h2f_ARLEN   : out   std_logic_vector(3 downto 0);                     -- arlen
			h2f_ARSIZE  : out   std_logic_vector(2 downto 0);                     -- arsize
			h2f_ARBURST : out   std_logic_vector(1 downto 0);                     -- arburst
			h2f_ARLOCK  : out   std_logic_vector(1 downto 0);                     -- arlock
			h2f_ARCACHE : out   std_logic_vector(3 downto 0);                     -- arcache
			h2f_ARPROT  : out   std_logic_vector(2 downto 0);                     -- arprot
			h2f_ARVALID : out   std_logic;                                        -- arvalid
			h2f_ARREADY : in    std_logic                     := 'X';             -- arready
			h2f_RID     : in    std_logic_vector(11 downto 0) := (others => 'X'); -- rid
			h2f_RDATA   : in    std_logic_vector(31 downto 0) := (others => 'X'); -- rdata
			h2f_RRESP   : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			h2f_RLAST   : in    std_logic                     := 'X';             -- rlast
			h2f_RVALID  : in    std_logic                     := 'X';             -- rvalid
			h2f_RREADY  : out   std_logic                                         -- rready
		);
	end component jaxa_hps_0;

	component jaxa_linkStatus is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(15 downto 0) := (others => 'X')  -- export
		);
	end component jaxa_linkStatus;

	component jaxa_pll_0 is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component jaxa_pll_0;

	component jaxa_receiveActivity is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic                     := 'X'              -- export
		);
	end component jaxa_receiveActivity;

	component jaxa_receiveFIFODataOut is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(8 downto 0)  := (others => 'X')  -- export
		);
	end component jaxa_receiveFIFODataOut;

	component jaxa_statisticalInformation_0 is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(31 downto 0) := (others => 'X')  -- export
		);
	end component jaxa_statisticalInformation_0;

	component jaxa_timeIn is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(5 downto 0)                      -- export
		);
	end component jaxa_timeIn;

	component jaxa_transmitFIFODataIn is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(8 downto 0)                      -- export
		);
	end component jaxa_transmitFIFODataIn;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal hps_0_h2f_reset_reset                    : std_logic; -- hps_0:h2f_rst_n -> hps_0_h2f_reset_reset:in
	signal rst_controller_reset_out_reset           : std_logic; -- rst_controller:reset_out -> rst_controller_reset_out_reset:in
	signal hps_0_h2f_reset_reset_ports_inv          : std_logic; -- hps_0_h2f_reset_reset:inv -> [pll_0:rst, rst_controller:reset_in0]
	signal rst_controller_reset_out_reset_ports_inv : std_logic; -- rst_controller_reset_out_reset:inv -> [autoStart:reset_n, controlFlagsIn:reset_n, controlFlagsOut:reset_n, creditCount:reset_n, errorStatus:reset_n, linkDisable:reset_n, linkStart:reset_n, linkStatus:reset_n, outstandingCount:reset_n, receiveActivity:reset_n, receiveClock:reset_n, receiveFIFODataCount:reset_n, receiveFIFODataOut:reset_n, receiveFIFOEmpty:reset_n, receiveFIFOFull:reset_n, receiveFIFOReadEnable:reset_n, spaceWireDataIn:reset_n, spaceWireDataOut:reset_n, spaceWireStrobeIn:reset_n, spaceWireStrobeOut:reset_n, statisticalInformationClear:reset_n, statisticalInformation_0:reset_n, statisticalInformation_1:reset_n, statisticalInformation_2:reset_n, statisticalInformation_3:reset_n, statisticalInformation_4:reset_n, statisticalInformation_5:reset_n, statisticalInformation_6:reset_n, statisticalInformation_7:reset_n, tickIn:reset_n, tickOut:reset_n, timeIn:reset_n, timeOut:reset_n, transmitActivity:reset_n, transmitClock:reset_n, transmitClockDivideValue:reset_n, transmitFIFODataCount:reset_n, transmitFIFODataIn:reset_n, transmitFIFOFull:reset_n, transmitFIFOWriteEnable:reset_n]

begin

	autostart : component jaxa_autoStart
		port map (
			clk        => clk_clk,                                  --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address    => open,                                     --                  s1.address
			write_n    => open,                                     --                    .write_n
			writedata  => open,                                     --                    .writedata
			chipselect => open,                                     --                    .chipselect
			readdata   => open,                                     --                    .readdata
			out_port   => autostart_external_connection_export      -- external_connection.export
		);

	controlflagsin : component jaxa_controlFlagsIn
		port map (
			clk        => clk_clk,                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => open,                                      --                  s1.address
			write_n    => open,                                      --                    .write_n
			writedata  => open,                                      --                    .writedata
			chipselect => open,                                      --                    .chipselect
			readdata   => open,                                      --                    .readdata
			out_port   => controlflagsin_external_connection_export  -- external_connection.export
		);

	controlflagsout : component jaxa_controlFlagsOut
		port map (
			clk      => clk_clk,                                    --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address  => open,                                       --                  s1.address
			readdata => open,                                       --                    .readdata
			in_port  => controlflagsout_external_connection_export  -- external_connection.export
		);

	creditcount : component jaxa_creditCount
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => open,                                     --                  s1.address
			readdata => open,                                     --                    .readdata
			in_port  => creditcount_external_connection_export    -- external_connection.export
		);

	errorstatus : component jaxa_errorStatus
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => open,                                     --                  s1.address
			readdata => open,                                     --                    .readdata
			in_port  => errorstatus_external_connection_export    -- external_connection.export
		);

	hps_0 : component jaxa_hps_0
		generic map (
			F2S_Width => 0,
			S2F_Width => 1
		)
		port map (
			mem_a       => memory_mem_a,          --         memory.mem_a
			mem_ba      => memory_mem_ba,         --               .mem_ba
			mem_ck      => memory_mem_ck,         --               .mem_ck
			mem_ck_n    => memory_mem_ck_n,       --               .mem_ck_n
			mem_cke     => memory_mem_cke,        --               .mem_cke
			mem_cs_n    => memory_mem_cs_n,       --               .mem_cs_n
			mem_ras_n   => memory_mem_ras_n,      --               .mem_ras_n
			mem_cas_n   => memory_mem_cas_n,      --               .mem_cas_n
			mem_we_n    => memory_mem_we_n,       --               .mem_we_n
			mem_reset_n => memory_mem_reset_n,    --               .mem_reset_n
			mem_dq      => memory_mem_dq,         --               .mem_dq
			mem_dqs     => memory_mem_dqs,        --               .mem_dqs
			mem_dqs_n   => memory_mem_dqs_n,      --               .mem_dqs_n
			mem_odt     => memory_mem_odt,        --               .mem_odt
			mem_dm      => memory_mem_dm,         --               .mem_dm
			oct_rzqin   => memory_oct_rzqin,      --               .oct_rzqin
			h2f_rst_n   => hps_0_h2f_reset_reset, --      h2f_reset.reset_n
			h2f_axi_clk => clk_clk,               --  h2f_axi_clock.clk
			h2f_AWID    => open,                  -- h2f_axi_master.awid
			h2f_AWADDR  => open,                  --               .awaddr
			h2f_AWLEN   => open,                  --               .awlen
			h2f_AWSIZE  => open,                  --               .awsize
			h2f_AWBURST => open,                  --               .awburst
			h2f_AWLOCK  => open,                  --               .awlock
			h2f_AWCACHE => open,                  --               .awcache
			h2f_AWPROT  => open,                  --               .awprot
			h2f_AWVALID => open,                  --               .awvalid
			h2f_AWREADY => open,                  --               .awready
			h2f_WID     => open,                  --               .wid
			h2f_WDATA   => open,                  --               .wdata
			h2f_WSTRB   => open,                  --               .wstrb
			h2f_WLAST   => open,                  --               .wlast
			h2f_WVALID  => open,                  --               .wvalid
			h2f_WREADY  => open,                  --               .wready
			h2f_BID     => open,                  --               .bid
			h2f_BRESP   => open,                  --               .bresp
			h2f_BVALID  => open,                  --               .bvalid
			h2f_BREADY  => open,                  --               .bready
			h2f_ARID    => open,                  --               .arid
			h2f_ARADDR  => open,                  --               .araddr
			h2f_ARLEN   => open,                  --               .arlen
			h2f_ARSIZE  => open,                  --               .arsize
			h2f_ARBURST => open,                  --               .arburst
			h2f_ARLOCK  => open,                  --               .arlock
			h2f_ARCACHE => open,                  --               .arcache
			h2f_ARPROT  => open,                  --               .arprot
			h2f_ARVALID => open,                  --               .arvalid
			h2f_ARREADY => open,                  --               .arready
			h2f_RID     => open,                  --               .rid
			h2f_RDATA   => open,                  --               .rdata
			h2f_RRESP   => open,                  --               .rresp
			h2f_RLAST   => open,                  --               .rlast
			h2f_RVALID  => open,                  --               .rvalid
			h2f_RREADY  => open                   --               .rready
		);

	linkdisable : component jaxa_autoStart
		port map (
			clk        => clk_clk,                                  --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address    => open,                                     --                  s1.address
			write_n    => open,                                     --                    .write_n
			writedata  => open,                                     --                    .writedata
			chipselect => open,                                     --                    .chipselect
			readdata   => open,                                     --                    .readdata
			out_port   => linkdisable_external_connection_export    -- external_connection.export
		);

	linkstart : component jaxa_autoStart
		port map (
			clk        => clk_clk,                                  --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address    => open,                                     --                  s1.address
			write_n    => open,                                     --                    .write_n
			writedata  => open,                                     --                    .writedata
			chipselect => open,                                     --                    .chipselect
			readdata   => open,                                     --                    .readdata
			out_port   => linkstart_external_connection_export      -- external_connection.export
		);

	linkstatus : component jaxa_linkStatus
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => open,                                     --                  s1.address
			readdata => open,                                     --                    .readdata
			in_port  => linkstatus_external_connection_export     -- external_connection.export
		);

	outstandingcount : component jaxa_creditCount
		port map (
			clk      => clk_clk,                                     --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address  => open,                                        --                  s1.address
			readdata => open,                                        --                    .readdata
			in_port  => outstandingcount_external_connection_export  -- external_connection.export
		);

	pll_0 : component jaxa_pll_0
		port map (
			refclk   => clk_clk,                         --  refclk.clk
			rst      => hps_0_h2f_reset_reset_ports_inv, --   reset.reset
			outclk_0 => pll_0_outclk0_clk,               -- outclk0.clk
			locked   => open                             --  locked.export
		);

	receiveactivity : component jaxa_receiveActivity
		port map (
			clk      => clk_clk,                                    --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address  => open,                                       --                  s1.address
			readdata => open,                                       --                    .readdata
			in_port  => receiveactivity_external_connection_export  -- external_connection.export
		);

	receiveclock : component jaxa_autoStart
		port map (
			clk        => clk_clk,                                  --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address    => open,                                     --                  s1.address
			write_n    => open,                                     --                    .write_n
			writedata  => open,                                     --                    .writedata
			chipselect => open,                                     --                    .chipselect
			readdata   => open,                                     --                    .readdata
			out_port   => receiveclock_external_connection_export   -- external_connection.export
		);

	receivefifodatacount : component jaxa_receiveActivity
		port map (
			clk      => clk_clk,                                         --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,        --               reset.reset_n
			address  => open,                                            --                  s1.address
			readdata => open,                                            --                    .readdata
			in_port  => receivefifodatacount_external_connection_export  -- external_connection.export
		);

	receivefifodataout : component jaxa_receiveFIFODataOut
		port map (
			clk      => clk_clk,                                       --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,      --               reset.reset_n
			address  => open,                                          --                  s1.address
			readdata => open,                                          --                    .readdata
			in_port  => receivefifodataout_external_connection_export  -- external_connection.export
		);

	receivefifoempty : component jaxa_receiveActivity
		port map (
			clk      => clk_clk,                                     --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address  => open,                                        --                  s1.address
			readdata => open,                                        --                    .readdata
			in_port  => receivefifoempty_external_connection_export  -- external_connection.export
		);

	receivefifofull : component jaxa_receiveActivity
		port map (
			clk      => clk_clk,                                    --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address  => open,                                       --                  s1.address
			readdata => open,                                       --                    .readdata
			in_port  => receivefifofull_external_connection_export  -- external_connection.export
		);

	receivefiforeadenable : component jaxa_autoStart
		port map (
			clk        => clk_clk,                                          --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,         --               reset.reset_n
			address    => open,                                             --                  s1.address
			write_n    => open,                                             --                    .write_n
			writedata  => open,                                             --                    .writedata
			chipselect => open,                                             --                    .chipselect
			readdata   => open,                                             --                    .readdata
			out_port   => receivefiforeadenable_external_connection_export  -- external_connection.export
		);

	spacewiredatain : component jaxa_autoStart
		port map (
			clk        => clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => open,                                       --                  s1.address
			write_n    => open,                                       --                    .write_n
			writedata  => open,                                       --                    .writedata
			chipselect => open,                                       --                    .chipselect
			readdata   => open,                                       --                    .readdata
			out_port   => spacewiredatain_external_connection_export  -- external_connection.export
		);

	spacewiredataout : component jaxa_receiveActivity
		port map (
			clk      => clk_clk,                                     --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address  => open,                                        --                  s1.address
			readdata => open,                                        --                    .readdata
			in_port  => spacewiredataout_external_connection_export  -- external_connection.export
		);

	spacewirestrobein : component jaxa_autoStart
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => open,                                         --                  s1.address
			write_n    => open,                                         --                    .write_n
			writedata  => open,                                         --                    .writedata
			chipselect => open,                                         --                    .chipselect
			readdata   => open,                                         --                    .readdata
			out_port   => spacewirestrobein_external_connection_export  -- external_connection.export
		);

	spacewirestrobeout : component jaxa_receiveActivity
		port map (
			clk      => clk_clk,                                       --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,      --               reset.reset_n
			address  => open,                                          --                  s1.address
			readdata => open,                                          --                    .readdata
			in_port  => spacewirestrobeout_external_connection_export  -- external_connection.export
		);

	statisticalinformationclear : component jaxa_autoStart
		port map (
			clk        => clk_clk,                                                --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,               --               reset.reset_n
			address    => open,                                                   --                  s1.address
			write_n    => open,                                                   --                    .write_n
			writedata  => open,                                                   --                    .writedata
			chipselect => open,                                                   --                    .chipselect
			readdata   => open,                                                   --                    .readdata
			out_port   => statisticalinformationclear_external_connection_export  -- external_connection.export
		);

	statisticalinformation_0 : component jaxa_statisticalInformation_0
		port map (
			clk      => clk_clk,                                             --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,            --               reset.reset_n
			address  => open,                                                --                  s1.address
			readdata => open,                                                --                    .readdata
			in_port  => statisticalinformation_0_external_connection_export  -- external_connection.export
		);

	statisticalinformation_1 : component jaxa_statisticalInformation_0
		port map (
			clk      => clk_clk,                                             --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,            --               reset.reset_n
			address  => open,                                                --                  s1.address
			readdata => open,                                                --                    .readdata
			in_port  => statisticalinformation_1_external_connection_export  -- external_connection.export
		);

	statisticalinformation_2 : component jaxa_statisticalInformation_0
		port map (
			clk      => clk_clk,                                             --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,            --               reset.reset_n
			address  => open,                                                --                  s1.address
			readdata => open,                                                --                    .readdata
			in_port  => statisticalinformation_2_external_connection_export  -- external_connection.export
		);

	statisticalinformation_3 : component jaxa_statisticalInformation_0
		port map (
			clk      => clk_clk,                                             --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,            --               reset.reset_n
			address  => open,                                                --                  s1.address
			readdata => open,                                                --                    .readdata
			in_port  => statisticalinformation_3_external_connection_export  -- external_connection.export
		);

	statisticalinformation_4 : component jaxa_statisticalInformation_0
		port map (
			clk      => clk_clk,                                             --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,            --               reset.reset_n
			address  => open,                                                --                  s1.address
			readdata => open,                                                --                    .readdata
			in_port  => statisticalinformation_4_external_connection_export  -- external_connection.export
		);

	statisticalinformation_5 : component jaxa_statisticalInformation_0
		port map (
			clk      => clk_clk,                                             --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,            --               reset.reset_n
			address  => open,                                                --                  s1.address
			readdata => open,                                                --                    .readdata
			in_port  => statisticalinformation_5_external_connection_export  -- external_connection.export
		);

	statisticalinformation_6 : component jaxa_statisticalInformation_0
		port map (
			clk      => clk_clk,                                             --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,            --               reset.reset_n
			address  => open,                                                --                  s1.address
			readdata => open,                                                --                    .readdata
			in_port  => statisticalinformation_6_external_connection_export  -- external_connection.export
		);

	statisticalinformation_7 : component jaxa_statisticalInformation_0
		port map (
			clk      => clk_clk,                                             --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,            --               reset.reset_n
			address  => open,                                                --                  s1.address
			readdata => open,                                                --                    .readdata
			in_port  => statisticalinformation_7_external_connection_export  -- external_connection.export
		);

	tickin : component jaxa_autoStart
		port map (
			clk        => clk_clk,                                  --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address    => open,                                     --                  s1.address
			write_n    => open,                                     --                    .write_n
			writedata  => open,                                     --                    .writedata
			chipselect => open,                                     --                    .chipselect
			readdata   => open,                                     --                    .readdata
			out_port   => tickin_external_connection_export         -- external_connection.export
		);

	tickout : component jaxa_receiveActivity
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => open,                                     --                  s1.address
			readdata => open,                                     --                    .readdata
			in_port  => tickout_external_connection_export        -- external_connection.export
		);

	timein : component jaxa_timeIn
		port map (
			clk        => clk_clk,                                  --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address    => open,                                     --                  s1.address
			write_n    => open,                                     --                    .write_n
			writedata  => open,                                     --                    .writedata
			chipselect => open,                                     --                    .chipselect
			readdata   => open,                                     --                    .readdata
			out_port   => timein_external_connection_export         -- external_connection.export
		);

	timeout : component jaxa_creditCount
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => open,                                     --                  s1.address
			readdata => open,                                     --                    .readdata
			in_port  => timeout_external_connection_export        -- external_connection.export
		);

	transmitactivity : component jaxa_receiveActivity
		port map (
			clk      => clk_clk,                                     --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address  => open,                                        --                  s1.address
			readdata => open,                                        --                    .readdata
			in_port  => transmitactivity_external_connection_export  -- external_connection.export
		);

	transmitclock : component jaxa_autoStart
		port map (
			clk        => clk_clk,                                  --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address    => open,                                     --                  s1.address
			write_n    => open,                                     --                    .write_n
			writedata  => open,                                     --                    .writedata
			chipselect => open,                                     --                    .chipselect
			readdata   => open,                                     --                    .readdata
			out_port   => transmitclock_external_connection_export  -- external_connection.export
		);

	transmitclockdividevalue : component jaxa_timeIn
		port map (
			clk        => clk_clk,                                             --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,            --               reset.reset_n
			address    => open,                                                --                  s1.address
			write_n    => open,                                                --                    .write_n
			writedata  => open,                                                --                    .writedata
			chipselect => open,                                                --                    .chipselect
			readdata   => open,                                                --                    .readdata
			out_port   => transmitclockdividevalue_external_connection_export  -- external_connection.export
		);

	transmitfifodatacount : component jaxa_creditCount
		port map (
			clk      => clk_clk,                                          --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,         --               reset.reset_n
			address  => open,                                             --                  s1.address
			readdata => open,                                             --                    .readdata
			in_port  => transmitfifodatacount_external_connection_export  -- external_connection.export
		);

	transmitfifodatain : component jaxa_transmitFIFODataIn
		port map (
			clk        => clk_clk,                                       --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,      --               reset.reset_n
			address    => open,                                          --                  s1.address
			write_n    => open,                                          --                    .write_n
			writedata  => open,                                          --                    .writedata
			chipselect => open,                                          --                    .chipselect
			readdata   => open,                                          --                    .readdata
			out_port   => transmitfifodatain_external_connection_export  -- external_connection.export
		);

	transmitfifofull : component jaxa_receiveActivity
		port map (
			clk      => clk_clk,                                     --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address  => open,                                        --                  s1.address
			readdata => open,                                        --                    .readdata
			in_port  => transmitfifofull_external_connection_export  -- external_connection.export
		);

	transmitfifowriteenable : component jaxa_autoStart
		port map (
			clk        => clk_clk,                                            --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,           --               reset.reset_n
			address    => open,                                               --                  s1.address
			write_n    => open,                                               --                    .write_n
			writedata  => open,                                               --                    .writedata
			chipselect => open,                                               --                    .chipselect
			readdata   => open,                                               --                    .readdata
			out_port   => transmitfifowriteenable_external_connection_export  -- external_connection.export
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => hps_0_h2f_reset_reset_ports_inv, -- reset_in0.reset
			clk            => clk_clk,                         --       clk.clk
			reset_out      => rst_controller_reset_out_reset,  -- reset_out.reset
			reset_req      => open,                            -- (terminated)
			reset_req_in0  => '0',                             -- (terminated)
			reset_in1      => '0',                             -- (terminated)
			reset_req_in1  => '0',                             -- (terminated)
			reset_in2      => '0',                             -- (terminated)
			reset_req_in2  => '0',                             -- (terminated)
			reset_in3      => '0',                             -- (terminated)
			reset_req_in3  => '0',                             -- (terminated)
			reset_in4      => '0',                             -- (terminated)
			reset_req_in4  => '0',                             -- (terminated)
			reset_in5      => '0',                             -- (terminated)
			reset_req_in5  => '0',                             -- (terminated)
			reset_in6      => '0',                             -- (terminated)
			reset_req_in6  => '0',                             -- (terminated)
			reset_in7      => '0',                             -- (terminated)
			reset_req_in7  => '0',                             -- (terminated)
			reset_in8      => '0',                             -- (terminated)
			reset_req_in8  => '0',                             -- (terminated)
			reset_in9      => '0',                             -- (terminated)
			reset_req_in9  => '0',                             -- (terminated)
			reset_in10     => '0',                             -- (terminated)
			reset_req_in10 => '0',                             -- (terminated)
			reset_in11     => '0',                             -- (terminated)
			reset_req_in11 => '0',                             -- (terminated)
			reset_in12     => '0',                             -- (terminated)
			reset_req_in12 => '0',                             -- (terminated)
			reset_in13     => '0',                             -- (terminated)
			reset_req_in13 => '0',                             -- (terminated)
			reset_in14     => '0',                             -- (terminated)
			reset_req_in14 => '0',                             -- (terminated)
			reset_in15     => '0',                             -- (terminated)
			reset_req_in15 => '0'                              -- (terminated)
		);

	hps_0_h2f_reset_reset_ports_inv <= not hps_0_h2f_reset_reset;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of jaxa
