// spw_babasu.v

// Generated using ACDS version 17.1 593

`timescale 1 ps / 1 ps
module spw_babasu (
		output wire        autostart_external_connection_export,    //    autostart_external_connection.export
		input  wire        clk_clk,                                 //                              clk.clk
		input  wire [2:0]  currentstate_external_connection_export, // currentstate_external_connection.export
		output wire [8:0]  data_i_external_connection_export,       //       data_i_external_connection.export
		input  wire [8:0]  data_o_external_connection_export,       //       data_o_external_connection.export
		input  wire [10:0] flags_external_connection_export,        //        flags_external_connection.export
		output wire        link_disable_external_connection_export, // link_disable_external_connection.export
		output wire        link_start_external_connection_export,   //   link_start_external_connection.export
		output wire        pll_0_outclk0_clk,                       //                    pll_0_outclk0.clk
		output wire        rd_data_external_connection_export,      //      rd_data_external_connection.export
		input  wire        reset_reset_n,                           //                            reset.reset_n
		input  wire        rx_empty_external_connection_export,     //     rx_empty_external_connection.export
		output wire        spill_enable_external_connection_export, // spill_enable_external_connection.export
		output wire        tick_in_external_connection_export,      //      tick_in_external_connection.export
		input  wire        tick_out_external_connection_export,     //     tick_out_external_connection.export
		output wire [7:0]  time_in_external_connection_export,      //      time_in_external_connection.export
		input  wire [7:0]  time_out_external_connection_export,     //     time_out_external_connection.export
		output wire [6:0]  tx_clk_div_external_connection_export,   //   tx_clk_div_external_connection.export
		input  wire        tx_full_external_connection_export,      //      tx_full_external_connection.export
		output wire        wr_data_external_connection_export       //      wr_data_external_connection.export
	);

	wire   [1:0] hps_0_h2f_axi_master_awburst;                 // hps_0:h2f_AWBURST -> mm_interconnect_0:hps_0_h2f_axi_master_awburst
	wire   [3:0] hps_0_h2f_axi_master_arlen;                   // hps_0:h2f_ARLEN -> mm_interconnect_0:hps_0_h2f_axi_master_arlen
	wire   [3:0] hps_0_h2f_axi_master_wstrb;                   // hps_0:h2f_WSTRB -> mm_interconnect_0:hps_0_h2f_axi_master_wstrb
	wire         hps_0_h2f_axi_master_wready;                  // mm_interconnect_0:hps_0_h2f_axi_master_wready -> hps_0:h2f_WREADY
	wire  [11:0] hps_0_h2f_axi_master_rid;                     // mm_interconnect_0:hps_0_h2f_axi_master_rid -> hps_0:h2f_RID
	wire         hps_0_h2f_axi_master_rready;                  // hps_0:h2f_RREADY -> mm_interconnect_0:hps_0_h2f_axi_master_rready
	wire   [3:0] hps_0_h2f_axi_master_awlen;                   // hps_0:h2f_AWLEN -> mm_interconnect_0:hps_0_h2f_axi_master_awlen
	wire  [11:0] hps_0_h2f_axi_master_wid;                     // hps_0:h2f_WID -> mm_interconnect_0:hps_0_h2f_axi_master_wid
	wire   [3:0] hps_0_h2f_axi_master_arcache;                 // hps_0:h2f_ARCACHE -> mm_interconnect_0:hps_0_h2f_axi_master_arcache
	wire         hps_0_h2f_axi_master_wvalid;                  // hps_0:h2f_WVALID -> mm_interconnect_0:hps_0_h2f_axi_master_wvalid
	wire  [29:0] hps_0_h2f_axi_master_araddr;                  // hps_0:h2f_ARADDR -> mm_interconnect_0:hps_0_h2f_axi_master_araddr
	wire   [2:0] hps_0_h2f_axi_master_arprot;                  // hps_0:h2f_ARPROT -> mm_interconnect_0:hps_0_h2f_axi_master_arprot
	wire   [2:0] hps_0_h2f_axi_master_awprot;                  // hps_0:h2f_AWPROT -> mm_interconnect_0:hps_0_h2f_axi_master_awprot
	wire  [31:0] hps_0_h2f_axi_master_wdata;                   // hps_0:h2f_WDATA -> mm_interconnect_0:hps_0_h2f_axi_master_wdata
	wire         hps_0_h2f_axi_master_arvalid;                 // hps_0:h2f_ARVALID -> mm_interconnect_0:hps_0_h2f_axi_master_arvalid
	wire   [3:0] hps_0_h2f_axi_master_awcache;                 // hps_0:h2f_AWCACHE -> mm_interconnect_0:hps_0_h2f_axi_master_awcache
	wire  [11:0] hps_0_h2f_axi_master_arid;                    // hps_0:h2f_ARID -> mm_interconnect_0:hps_0_h2f_axi_master_arid
	wire   [1:0] hps_0_h2f_axi_master_arlock;                  // hps_0:h2f_ARLOCK -> mm_interconnect_0:hps_0_h2f_axi_master_arlock
	wire   [1:0] hps_0_h2f_axi_master_awlock;                  // hps_0:h2f_AWLOCK -> mm_interconnect_0:hps_0_h2f_axi_master_awlock
	wire  [29:0] hps_0_h2f_axi_master_awaddr;                  // hps_0:h2f_AWADDR -> mm_interconnect_0:hps_0_h2f_axi_master_awaddr
	wire   [1:0] hps_0_h2f_axi_master_bresp;                   // mm_interconnect_0:hps_0_h2f_axi_master_bresp -> hps_0:h2f_BRESP
	wire         hps_0_h2f_axi_master_arready;                 // mm_interconnect_0:hps_0_h2f_axi_master_arready -> hps_0:h2f_ARREADY
	wire  [31:0] hps_0_h2f_axi_master_rdata;                   // mm_interconnect_0:hps_0_h2f_axi_master_rdata -> hps_0:h2f_RDATA
	wire         hps_0_h2f_axi_master_awready;                 // mm_interconnect_0:hps_0_h2f_axi_master_awready -> hps_0:h2f_AWREADY
	wire   [1:0] hps_0_h2f_axi_master_arburst;                 // hps_0:h2f_ARBURST -> mm_interconnect_0:hps_0_h2f_axi_master_arburst
	wire   [2:0] hps_0_h2f_axi_master_arsize;                  // hps_0:h2f_ARSIZE -> mm_interconnect_0:hps_0_h2f_axi_master_arsize
	wire         hps_0_h2f_axi_master_bready;                  // hps_0:h2f_BREADY -> mm_interconnect_0:hps_0_h2f_axi_master_bready
	wire         hps_0_h2f_axi_master_rlast;                   // mm_interconnect_0:hps_0_h2f_axi_master_rlast -> hps_0:h2f_RLAST
	wire         hps_0_h2f_axi_master_wlast;                   // hps_0:h2f_WLAST -> mm_interconnect_0:hps_0_h2f_axi_master_wlast
	wire   [1:0] hps_0_h2f_axi_master_rresp;                   // mm_interconnect_0:hps_0_h2f_axi_master_rresp -> hps_0:h2f_RRESP
	wire  [11:0] hps_0_h2f_axi_master_awid;                    // hps_0:h2f_AWID -> mm_interconnect_0:hps_0_h2f_axi_master_awid
	wire  [11:0] hps_0_h2f_axi_master_bid;                     // mm_interconnect_0:hps_0_h2f_axi_master_bid -> hps_0:h2f_BID
	wire         hps_0_h2f_axi_master_bvalid;                  // mm_interconnect_0:hps_0_h2f_axi_master_bvalid -> hps_0:h2f_BVALID
	wire   [2:0] hps_0_h2f_axi_master_awsize;                  // hps_0:h2f_AWSIZE -> mm_interconnect_0:hps_0_h2f_axi_master_awsize
	wire         hps_0_h2f_axi_master_awvalid;                 // hps_0:h2f_AWVALID -> mm_interconnect_0:hps_0_h2f_axi_master_awvalid
	wire         hps_0_h2f_axi_master_rvalid;                  // mm_interconnect_0:hps_0_h2f_axi_master_rvalid -> hps_0:h2f_RVALID
	wire         mm_interconnect_0_link_start_s1_chipselect;   // mm_interconnect_0:LINK_START_s1_chipselect -> LINK_START:chipselect
	wire  [31:0] mm_interconnect_0_link_start_s1_readdata;     // LINK_START:readdata -> mm_interconnect_0:LINK_START_s1_readdata
	wire   [1:0] mm_interconnect_0_link_start_s1_address;      // mm_interconnect_0:LINK_START_s1_address -> LINK_START:address
	wire         mm_interconnect_0_link_start_s1_write;        // mm_interconnect_0:LINK_START_s1_write -> LINK_START:write_n
	wire  [31:0] mm_interconnect_0_link_start_s1_writedata;    // mm_interconnect_0:LINK_START_s1_writedata -> LINK_START:writedata
	wire         mm_interconnect_0_link_disable_s1_chipselect; // mm_interconnect_0:LINK_DISABLE_s1_chipselect -> LINK_DISABLE:chipselect
	wire  [31:0] mm_interconnect_0_link_disable_s1_readdata;   // LINK_DISABLE:readdata -> mm_interconnect_0:LINK_DISABLE_s1_readdata
	wire   [1:0] mm_interconnect_0_link_disable_s1_address;    // mm_interconnect_0:LINK_DISABLE_s1_address -> LINK_DISABLE:address
	wire         mm_interconnect_0_link_disable_s1_write;      // mm_interconnect_0:LINK_DISABLE_s1_write -> LINK_DISABLE:write_n
	wire  [31:0] mm_interconnect_0_link_disable_s1_writedata;  // mm_interconnect_0:LINK_DISABLE_s1_writedata -> LINK_DISABLE:writedata
	wire         mm_interconnect_0_autostart_s1_chipselect;    // mm_interconnect_0:AUTOSTART_s1_chipselect -> AUTOSTART:chipselect
	wire  [31:0] mm_interconnect_0_autostart_s1_readdata;      // AUTOSTART:readdata -> mm_interconnect_0:AUTOSTART_s1_readdata
	wire   [1:0] mm_interconnect_0_autostart_s1_address;       // mm_interconnect_0:AUTOSTART_s1_address -> AUTOSTART:address
	wire         mm_interconnect_0_autostart_s1_write;         // mm_interconnect_0:AUTOSTART_s1_write -> AUTOSTART:write_n
	wire  [31:0] mm_interconnect_0_autostart_s1_writedata;     // mm_interconnect_0:AUTOSTART_s1_writedata -> AUTOSTART:writedata
	wire  [31:0] mm_interconnect_0_currentstate_s1_readdata;   // CURRENTSTATE:readdata -> mm_interconnect_0:CURRENTSTATE_s1_readdata
	wire   [1:0] mm_interconnect_0_currentstate_s1_address;    // mm_interconnect_0:CURRENTSTATE_s1_address -> CURRENTSTATE:address
	wire  [31:0] mm_interconnect_0_flags_s1_readdata;          // FLAGS:readdata -> mm_interconnect_0:FLAGS_s1_readdata
	wire   [1:0] mm_interconnect_0_flags_s1_address;           // mm_interconnect_0:FLAGS_s1_address -> FLAGS:address
	wire         mm_interconnect_0_data_i_s1_chipselect;       // mm_interconnect_0:DATA_I_s1_chipselect -> DATA_I:chipselect
	wire  [31:0] mm_interconnect_0_data_i_s1_readdata;         // DATA_I:readdata -> mm_interconnect_0:DATA_I_s1_readdata
	wire   [1:0] mm_interconnect_0_data_i_s1_address;          // mm_interconnect_0:DATA_I_s1_address -> DATA_I:address
	wire         mm_interconnect_0_data_i_s1_write;            // mm_interconnect_0:DATA_I_s1_write -> DATA_I:write_n
	wire  [31:0] mm_interconnect_0_data_i_s1_writedata;        // mm_interconnect_0:DATA_I_s1_writedata -> DATA_I:writedata
	wire         mm_interconnect_0_wr_data_s1_chipselect;      // mm_interconnect_0:WR_DATA_s1_chipselect -> WR_DATA:chipselect
	wire  [31:0] mm_interconnect_0_wr_data_s1_readdata;        // WR_DATA:readdata -> mm_interconnect_0:WR_DATA_s1_readdata
	wire   [1:0] mm_interconnect_0_wr_data_s1_address;         // mm_interconnect_0:WR_DATA_s1_address -> WR_DATA:address
	wire         mm_interconnect_0_wr_data_s1_write;           // mm_interconnect_0:WR_DATA_s1_write -> WR_DATA:write_n
	wire  [31:0] mm_interconnect_0_wr_data_s1_writedata;       // mm_interconnect_0:WR_DATA_s1_writedata -> WR_DATA:writedata
	wire  [31:0] mm_interconnect_0_tx_full_s1_readdata;        // TX_FULL:readdata -> mm_interconnect_0:TX_FULL_s1_readdata
	wire   [1:0] mm_interconnect_0_tx_full_s1_address;         // mm_interconnect_0:TX_FULL_s1_address -> TX_FULL:address
	wire  [31:0] mm_interconnect_0_data_o_s1_readdata;         // DATA_O:readdata -> mm_interconnect_0:DATA_O_s1_readdata
	wire   [1:0] mm_interconnect_0_data_o_s1_address;          // mm_interconnect_0:DATA_O_s1_address -> DATA_O:address
	wire         mm_interconnect_0_rd_data_s1_chipselect;      // mm_interconnect_0:RD_DATA_s1_chipselect -> RD_DATA:chipselect
	wire  [31:0] mm_interconnect_0_rd_data_s1_readdata;        // RD_DATA:readdata -> mm_interconnect_0:RD_DATA_s1_readdata
	wire   [1:0] mm_interconnect_0_rd_data_s1_address;         // mm_interconnect_0:RD_DATA_s1_address -> RD_DATA:address
	wire         mm_interconnect_0_rd_data_s1_write;           // mm_interconnect_0:RD_DATA_s1_write -> RD_DATA:write_n
	wire  [31:0] mm_interconnect_0_rd_data_s1_writedata;       // mm_interconnect_0:RD_DATA_s1_writedata -> RD_DATA:writedata
	wire  [31:0] mm_interconnect_0_rx_empty_s1_readdata;       // RX_EMPTY:readdata -> mm_interconnect_0:RX_EMPTY_s1_readdata
	wire   [1:0] mm_interconnect_0_rx_empty_s1_address;        // mm_interconnect_0:RX_EMPTY_s1_address -> RX_EMPTY:address
	wire  [31:0] mm_interconnect_0_tick_out_s1_readdata;       // TICK_OUT:readdata -> mm_interconnect_0:TICK_OUT_s1_readdata
	wire   [1:0] mm_interconnect_0_tick_out_s1_address;        // mm_interconnect_0:TICK_OUT_s1_address -> TICK_OUT:address
	wire  [31:0] mm_interconnect_0_time_out_s1_readdata;       // TIME_OUT:readdata -> mm_interconnect_0:TIME_OUT_s1_readdata
	wire   [1:0] mm_interconnect_0_time_out_s1_address;        // mm_interconnect_0:TIME_OUT_s1_address -> TIME_OUT:address
	wire         mm_interconnect_0_tick_in_s1_chipselect;      // mm_interconnect_0:TICK_IN_s1_chipselect -> TICK_IN:chipselect
	wire  [31:0] mm_interconnect_0_tick_in_s1_readdata;        // TICK_IN:readdata -> mm_interconnect_0:TICK_IN_s1_readdata
	wire   [1:0] mm_interconnect_0_tick_in_s1_address;         // mm_interconnect_0:TICK_IN_s1_address -> TICK_IN:address
	wire         mm_interconnect_0_tick_in_s1_write;           // mm_interconnect_0:TICK_IN_s1_write -> TICK_IN:write_n
	wire  [31:0] mm_interconnect_0_tick_in_s1_writedata;       // mm_interconnect_0:TICK_IN_s1_writedata -> TICK_IN:writedata
	wire         mm_interconnect_0_time_in_s1_chipselect;      // mm_interconnect_0:TIME_IN_s1_chipselect -> TIME_IN:chipselect
	wire  [31:0] mm_interconnect_0_time_in_s1_readdata;        // TIME_IN:readdata -> mm_interconnect_0:TIME_IN_s1_readdata
	wire   [1:0] mm_interconnect_0_time_in_s1_address;         // mm_interconnect_0:TIME_IN_s1_address -> TIME_IN:address
	wire         mm_interconnect_0_time_in_s1_write;           // mm_interconnect_0:TIME_IN_s1_write -> TIME_IN:write_n
	wire  [31:0] mm_interconnect_0_time_in_s1_writedata;       // mm_interconnect_0:TIME_IN_s1_writedata -> TIME_IN:writedata
	wire         mm_interconnect_0_tx_clk_div_s1_chipselect;   // mm_interconnect_0:TX_CLK_DIV_s1_chipselect -> TX_CLK_DIV:chipselect
	wire  [31:0] mm_interconnect_0_tx_clk_div_s1_readdata;     // TX_CLK_DIV:readdata -> mm_interconnect_0:TX_CLK_DIV_s1_readdata
	wire   [1:0] mm_interconnect_0_tx_clk_div_s1_address;      // mm_interconnect_0:TX_CLK_DIV_s1_address -> TX_CLK_DIV:address
	wire         mm_interconnect_0_tx_clk_div_s1_write;        // mm_interconnect_0:TX_CLK_DIV_s1_write -> TX_CLK_DIV:write_n
	wire  [31:0] mm_interconnect_0_tx_clk_div_s1_writedata;    // mm_interconnect_0:TX_CLK_DIV_s1_writedata -> TX_CLK_DIV:writedata
	wire         mm_interconnect_0_spill_enable_s1_chipselect; // mm_interconnect_0:SPILL_ENABLE_s1_chipselect -> SPILL_ENABLE:chipselect
	wire  [31:0] mm_interconnect_0_spill_enable_s1_readdata;   // SPILL_ENABLE:readdata -> mm_interconnect_0:SPILL_ENABLE_s1_readdata
	wire   [1:0] mm_interconnect_0_spill_enable_s1_address;    // mm_interconnect_0:SPILL_ENABLE_s1_address -> SPILL_ENABLE:address
	wire         mm_interconnect_0_spill_enable_s1_write;      // mm_interconnect_0:SPILL_ENABLE_s1_write -> SPILL_ENABLE:write_n
	wire  [31:0] mm_interconnect_0_spill_enable_s1_writedata;  // mm_interconnect_0:SPILL_ENABLE_s1_writedata -> SPILL_ENABLE:writedata
	wire         rst_controller_reset_out_reset;               // rst_controller:reset_out -> [AUTOSTART:reset_n, CURRENTSTATE:reset_n, DATA_I:reset_n, DATA_O:reset_n, FLAGS:reset_n, LINK_DISABLE:reset_n, LINK_START:reset_n, RD_DATA:reset_n, RX_EMPTY:reset_n, SPILL_ENABLE:reset_n, TICK_IN:reset_n, TICK_OUT:reset_n, TIME_IN:reset_n, TIME_OUT:reset_n, TX_CLK_DIV:reset_n, TX_FULL:reset_n, WR_DATA:reset_n, mm_interconnect_0:LINK_START_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset;           // rst_controller_001:reset_out -> mm_interconnect_0:hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset
	wire         hps_0_h2f_reset_reset;                        // hps_0:h2f_rst_n -> rst_controller_001:reset_in0

	spw_babasu_AUTOSTART autostart (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_autostart_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_autostart_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_autostart_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_autostart_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_autostart_s1_readdata),   //                    .readdata
		.out_port   (autostart_external_connection_export)       // external_connection.export
	);

	spw_babasu_CURRENTSTATE currentstate (
		.clk      (clk_clk),                                    //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_0_currentstate_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_currentstate_s1_readdata), //                    .readdata
		.in_port  (currentstate_external_connection_export)     // external_connection.export
	);

	spw_babasu_DATA_I data_i (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_data_i_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_data_i_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_data_i_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_data_i_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_data_i_s1_readdata),   //                    .readdata
		.out_port   (data_i_external_connection_export)       // external_connection.export
	);

	spw_babasu_DATA_O data_o (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_data_o_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_data_o_s1_readdata), //                    .readdata
		.in_port  (data_o_external_connection_export)     // external_connection.export
	);

	spw_babasu_FLAGS flags (
		.clk      (clk_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_flags_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_flags_s1_readdata), //                    .readdata
		.in_port  (flags_external_connection_export)     // external_connection.export
	);

	spw_babasu_AUTOSTART link_disable (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_link_disable_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_link_disable_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_link_disable_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_link_disable_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_link_disable_s1_readdata),   //                    .readdata
		.out_port   (link_disable_external_connection_export)       // external_connection.export
	);

	spw_babasu_AUTOSTART link_start (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_link_start_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_link_start_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_link_start_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_link_start_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_link_start_s1_readdata),   //                    .readdata
		.out_port   (link_start_external_connection_export)       // external_connection.export
	);

	spw_babasu_AUTOSTART rd_data (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_rd_data_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_rd_data_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_rd_data_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_rd_data_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_rd_data_s1_readdata),   //                    .readdata
		.out_port   (rd_data_external_connection_export)       // external_connection.export
	);

	spw_babasu_RX_EMPTY rx_empty (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_rx_empty_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_rx_empty_s1_readdata), //                    .readdata
		.in_port  (rx_empty_external_connection_export)     // external_connection.export
	);

	spw_babasu_SPILL_ENABLE spill_enable (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_spill_enable_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_spill_enable_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_spill_enable_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_spill_enable_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_spill_enable_s1_readdata),   //                    .readdata
		.out_port   (spill_enable_external_connection_export)       // external_connection.export
	);

	spw_babasu_AUTOSTART tick_in (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_tick_in_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_tick_in_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_tick_in_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_tick_in_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_tick_in_s1_readdata),   //                    .readdata
		.out_port   (tick_in_external_connection_export)       // external_connection.export
	);

	spw_babasu_RX_EMPTY tick_out (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_tick_out_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_tick_out_s1_readdata), //                    .readdata
		.in_port  (tick_out_external_connection_export)     // external_connection.export
	);

	spw_babasu_TIME_IN time_in (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_time_in_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_time_in_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_time_in_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_time_in_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_time_in_s1_readdata),   //                    .readdata
		.out_port   (time_in_external_connection_export)       // external_connection.export
	);

	spw_babasu_TIME_OUT time_out (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_time_out_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_time_out_s1_readdata), //                    .readdata
		.in_port  (time_out_external_connection_export)     // external_connection.export
	);

	spw_babasu_TX_CLK_DIV tx_clk_div (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_tx_clk_div_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_tx_clk_div_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_tx_clk_div_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_tx_clk_div_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_tx_clk_div_s1_readdata),   //                    .readdata
		.out_port   (tx_clk_div_external_connection_export)       // external_connection.export
	);

	spw_babasu_RX_EMPTY tx_full (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_tx_full_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_tx_full_s1_readdata), //                    .readdata
		.in_port  (tx_full_external_connection_export)     // external_connection.export
	);

	spw_babasu_AUTOSTART wr_data (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_wr_data_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_wr_data_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_wr_data_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_wr_data_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_wr_data_s1_readdata),   //                    .readdata
		.out_port   (wr_data_external_connection_export)       // external_connection.export
	);

	spw_babasu_hps_0 #(
		.F2S_Width (0),
		.S2F_Width (1)
	) hps_0 (
		.mem_a       (),                             //         memory.mem_a
		.mem_ba      (),                             //               .mem_ba
		.mem_ck      (),                             //               .mem_ck
		.mem_ck_n    (),                             //               .mem_ck_n
		.mem_cke     (),                             //               .mem_cke
		.mem_cs_n    (),                             //               .mem_cs_n
		.mem_ras_n   (),                             //               .mem_ras_n
		.mem_cas_n   (),                             //               .mem_cas_n
		.mem_we_n    (),                             //               .mem_we_n
		.mem_reset_n (),                             //               .mem_reset_n
		.mem_dq      (),                             //               .mem_dq
		.mem_dqs     (),                             //               .mem_dqs
		.mem_dqs_n   (),                             //               .mem_dqs_n
		.mem_odt     (),                             //               .mem_odt
		.mem_dm      (),                             //               .mem_dm
		.oct_rzqin   (),                             //               .oct_rzqin
		.h2f_rst_n   (hps_0_h2f_reset_reset),        //      h2f_reset.reset_n
		.h2f_axi_clk (clk_clk),                      //  h2f_axi_clock.clk
		.h2f_AWID    (hps_0_h2f_axi_master_awid),    // h2f_axi_master.awid
		.h2f_AWADDR  (hps_0_h2f_axi_master_awaddr),  //               .awaddr
		.h2f_AWLEN   (hps_0_h2f_axi_master_awlen),   //               .awlen
		.h2f_AWSIZE  (hps_0_h2f_axi_master_awsize),  //               .awsize
		.h2f_AWBURST (hps_0_h2f_axi_master_awburst), //               .awburst
		.h2f_AWLOCK  (hps_0_h2f_axi_master_awlock),  //               .awlock
		.h2f_AWCACHE (hps_0_h2f_axi_master_awcache), //               .awcache
		.h2f_AWPROT  (hps_0_h2f_axi_master_awprot),  //               .awprot
		.h2f_AWVALID (hps_0_h2f_axi_master_awvalid), //               .awvalid
		.h2f_AWREADY (hps_0_h2f_axi_master_awready), //               .awready
		.h2f_WID     (hps_0_h2f_axi_master_wid),     //               .wid
		.h2f_WDATA   (hps_0_h2f_axi_master_wdata),   //               .wdata
		.h2f_WSTRB   (hps_0_h2f_axi_master_wstrb),   //               .wstrb
		.h2f_WLAST   (hps_0_h2f_axi_master_wlast),   //               .wlast
		.h2f_WVALID  (hps_0_h2f_axi_master_wvalid),  //               .wvalid
		.h2f_WREADY  (hps_0_h2f_axi_master_wready),  //               .wready
		.h2f_BID     (hps_0_h2f_axi_master_bid),     //               .bid
		.h2f_BRESP   (hps_0_h2f_axi_master_bresp),   //               .bresp
		.h2f_BVALID  (hps_0_h2f_axi_master_bvalid),  //               .bvalid
		.h2f_BREADY  (hps_0_h2f_axi_master_bready),  //               .bready
		.h2f_ARID    (hps_0_h2f_axi_master_arid),    //               .arid
		.h2f_ARADDR  (hps_0_h2f_axi_master_araddr),  //               .araddr
		.h2f_ARLEN   (hps_0_h2f_axi_master_arlen),   //               .arlen
		.h2f_ARSIZE  (hps_0_h2f_axi_master_arsize),  //               .arsize
		.h2f_ARBURST (hps_0_h2f_axi_master_arburst), //               .arburst
		.h2f_ARLOCK  (hps_0_h2f_axi_master_arlock),  //               .arlock
		.h2f_ARCACHE (hps_0_h2f_axi_master_arcache), //               .arcache
		.h2f_ARPROT  (hps_0_h2f_axi_master_arprot),  //               .arprot
		.h2f_ARVALID (hps_0_h2f_axi_master_arvalid), //               .arvalid
		.h2f_ARREADY (hps_0_h2f_axi_master_arready), //               .arready
		.h2f_RID     (hps_0_h2f_axi_master_rid),     //               .rid
		.h2f_RDATA   (hps_0_h2f_axi_master_rdata),   //               .rdata
		.h2f_RRESP   (hps_0_h2f_axi_master_rresp),   //               .rresp
		.h2f_RLAST   (hps_0_h2f_axi_master_rlast),   //               .rlast
		.h2f_RVALID  (hps_0_h2f_axi_master_rvalid),  //               .rvalid
		.h2f_RREADY  (hps_0_h2f_axi_master_rready)   //               .rready
	);

	spw_babasu_pll_0 pll_0 (
		.refclk   (clk_clk),           //  refclk.clk
		.rst      (~reset_reset_n),    //   reset.reset
		.outclk_0 (pll_0_outclk0_clk), // outclk0.clk
		.locked   ()                   // (terminated)
	);

	spw_babasu_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_h2f_axi_master_awid                                        (hps_0_h2f_axi_master_awid),                    //                                       hps_0_h2f_axi_master.awid
		.hps_0_h2f_axi_master_awaddr                                      (hps_0_h2f_axi_master_awaddr),                  //                                                           .awaddr
		.hps_0_h2f_axi_master_awlen                                       (hps_0_h2f_axi_master_awlen),                   //                                                           .awlen
		.hps_0_h2f_axi_master_awsize                                      (hps_0_h2f_axi_master_awsize),                  //                                                           .awsize
		.hps_0_h2f_axi_master_awburst                                     (hps_0_h2f_axi_master_awburst),                 //                                                           .awburst
		.hps_0_h2f_axi_master_awlock                                      (hps_0_h2f_axi_master_awlock),                  //                                                           .awlock
		.hps_0_h2f_axi_master_awcache                                     (hps_0_h2f_axi_master_awcache),                 //                                                           .awcache
		.hps_0_h2f_axi_master_awprot                                      (hps_0_h2f_axi_master_awprot),                  //                                                           .awprot
		.hps_0_h2f_axi_master_awvalid                                     (hps_0_h2f_axi_master_awvalid),                 //                                                           .awvalid
		.hps_0_h2f_axi_master_awready                                     (hps_0_h2f_axi_master_awready),                 //                                                           .awready
		.hps_0_h2f_axi_master_wid                                         (hps_0_h2f_axi_master_wid),                     //                                                           .wid
		.hps_0_h2f_axi_master_wdata                                       (hps_0_h2f_axi_master_wdata),                   //                                                           .wdata
		.hps_0_h2f_axi_master_wstrb                                       (hps_0_h2f_axi_master_wstrb),                   //                                                           .wstrb
		.hps_0_h2f_axi_master_wlast                                       (hps_0_h2f_axi_master_wlast),                   //                                                           .wlast
		.hps_0_h2f_axi_master_wvalid                                      (hps_0_h2f_axi_master_wvalid),                  //                                                           .wvalid
		.hps_0_h2f_axi_master_wready                                      (hps_0_h2f_axi_master_wready),                  //                                                           .wready
		.hps_0_h2f_axi_master_bid                                         (hps_0_h2f_axi_master_bid),                     //                                                           .bid
		.hps_0_h2f_axi_master_bresp                                       (hps_0_h2f_axi_master_bresp),                   //                                                           .bresp
		.hps_0_h2f_axi_master_bvalid                                      (hps_0_h2f_axi_master_bvalid),                  //                                                           .bvalid
		.hps_0_h2f_axi_master_bready                                      (hps_0_h2f_axi_master_bready),                  //                                                           .bready
		.hps_0_h2f_axi_master_arid                                        (hps_0_h2f_axi_master_arid),                    //                                                           .arid
		.hps_0_h2f_axi_master_araddr                                      (hps_0_h2f_axi_master_araddr),                  //                                                           .araddr
		.hps_0_h2f_axi_master_arlen                                       (hps_0_h2f_axi_master_arlen),                   //                                                           .arlen
		.hps_0_h2f_axi_master_arsize                                      (hps_0_h2f_axi_master_arsize),                  //                                                           .arsize
		.hps_0_h2f_axi_master_arburst                                     (hps_0_h2f_axi_master_arburst),                 //                                                           .arburst
		.hps_0_h2f_axi_master_arlock                                      (hps_0_h2f_axi_master_arlock),                  //                                                           .arlock
		.hps_0_h2f_axi_master_arcache                                     (hps_0_h2f_axi_master_arcache),                 //                                                           .arcache
		.hps_0_h2f_axi_master_arprot                                      (hps_0_h2f_axi_master_arprot),                  //                                                           .arprot
		.hps_0_h2f_axi_master_arvalid                                     (hps_0_h2f_axi_master_arvalid),                 //                                                           .arvalid
		.hps_0_h2f_axi_master_arready                                     (hps_0_h2f_axi_master_arready),                 //                                                           .arready
		.hps_0_h2f_axi_master_rid                                         (hps_0_h2f_axi_master_rid),                     //                                                           .rid
		.hps_0_h2f_axi_master_rdata                                       (hps_0_h2f_axi_master_rdata),                   //                                                           .rdata
		.hps_0_h2f_axi_master_rresp                                       (hps_0_h2f_axi_master_rresp),                   //                                                           .rresp
		.hps_0_h2f_axi_master_rlast                                       (hps_0_h2f_axi_master_rlast),                   //                                                           .rlast
		.hps_0_h2f_axi_master_rvalid                                      (hps_0_h2f_axi_master_rvalid),                  //                                                           .rvalid
		.hps_0_h2f_axi_master_rready                                      (hps_0_h2f_axi_master_rready),                  //                                                           .rready
		.clk_0_clk_clk                                                    (clk_clk),                                      //                                                  clk_0_clk.clk
		.hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),           // hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.LINK_START_reset_reset_bridge_in_reset_reset                     (rst_controller_reset_out_reset),               //                     LINK_START_reset_reset_bridge_in_reset.reset
		.AUTOSTART_s1_address                                             (mm_interconnect_0_autostart_s1_address),       //                                               AUTOSTART_s1.address
		.AUTOSTART_s1_write                                               (mm_interconnect_0_autostart_s1_write),         //                                                           .write
		.AUTOSTART_s1_readdata                                            (mm_interconnect_0_autostart_s1_readdata),      //                                                           .readdata
		.AUTOSTART_s1_writedata                                           (mm_interconnect_0_autostart_s1_writedata),     //                                                           .writedata
		.AUTOSTART_s1_chipselect                                          (mm_interconnect_0_autostart_s1_chipselect),    //                                                           .chipselect
		.CURRENTSTATE_s1_address                                          (mm_interconnect_0_currentstate_s1_address),    //                                            CURRENTSTATE_s1.address
		.CURRENTSTATE_s1_readdata                                         (mm_interconnect_0_currentstate_s1_readdata),   //                                                           .readdata
		.DATA_I_s1_address                                                (mm_interconnect_0_data_i_s1_address),          //                                                  DATA_I_s1.address
		.DATA_I_s1_write                                                  (mm_interconnect_0_data_i_s1_write),            //                                                           .write
		.DATA_I_s1_readdata                                               (mm_interconnect_0_data_i_s1_readdata),         //                                                           .readdata
		.DATA_I_s1_writedata                                              (mm_interconnect_0_data_i_s1_writedata),        //                                                           .writedata
		.DATA_I_s1_chipselect                                             (mm_interconnect_0_data_i_s1_chipselect),       //                                                           .chipselect
		.DATA_O_s1_address                                                (mm_interconnect_0_data_o_s1_address),          //                                                  DATA_O_s1.address
		.DATA_O_s1_readdata                                               (mm_interconnect_0_data_o_s1_readdata),         //                                                           .readdata
		.FLAGS_s1_address                                                 (mm_interconnect_0_flags_s1_address),           //                                                   FLAGS_s1.address
		.FLAGS_s1_readdata                                                (mm_interconnect_0_flags_s1_readdata),          //                                                           .readdata
		.LINK_DISABLE_s1_address                                          (mm_interconnect_0_link_disable_s1_address),    //                                            LINK_DISABLE_s1.address
		.LINK_DISABLE_s1_write                                            (mm_interconnect_0_link_disable_s1_write),      //                                                           .write
		.LINK_DISABLE_s1_readdata                                         (mm_interconnect_0_link_disable_s1_readdata),   //                                                           .readdata
		.LINK_DISABLE_s1_writedata                                        (mm_interconnect_0_link_disable_s1_writedata),  //                                                           .writedata
		.LINK_DISABLE_s1_chipselect                                       (mm_interconnect_0_link_disable_s1_chipselect), //                                                           .chipselect
		.LINK_START_s1_address                                            (mm_interconnect_0_link_start_s1_address),      //                                              LINK_START_s1.address
		.LINK_START_s1_write                                              (mm_interconnect_0_link_start_s1_write),        //                                                           .write
		.LINK_START_s1_readdata                                           (mm_interconnect_0_link_start_s1_readdata),     //                                                           .readdata
		.LINK_START_s1_writedata                                          (mm_interconnect_0_link_start_s1_writedata),    //                                                           .writedata
		.LINK_START_s1_chipselect                                         (mm_interconnect_0_link_start_s1_chipselect),   //                                                           .chipselect
		.RD_DATA_s1_address                                               (mm_interconnect_0_rd_data_s1_address),         //                                                 RD_DATA_s1.address
		.RD_DATA_s1_write                                                 (mm_interconnect_0_rd_data_s1_write),           //                                                           .write
		.RD_DATA_s1_readdata                                              (mm_interconnect_0_rd_data_s1_readdata),        //                                                           .readdata
		.RD_DATA_s1_writedata                                             (mm_interconnect_0_rd_data_s1_writedata),       //                                                           .writedata
		.RD_DATA_s1_chipselect                                            (mm_interconnect_0_rd_data_s1_chipselect),      //                                                           .chipselect
		.RX_EMPTY_s1_address                                              (mm_interconnect_0_rx_empty_s1_address),        //                                                RX_EMPTY_s1.address
		.RX_EMPTY_s1_readdata                                             (mm_interconnect_0_rx_empty_s1_readdata),       //                                                           .readdata
		.SPILL_ENABLE_s1_address                                          (mm_interconnect_0_spill_enable_s1_address),    //                                            SPILL_ENABLE_s1.address
		.SPILL_ENABLE_s1_write                                            (mm_interconnect_0_spill_enable_s1_write),      //                                                           .write
		.SPILL_ENABLE_s1_readdata                                         (mm_interconnect_0_spill_enable_s1_readdata),   //                                                           .readdata
		.SPILL_ENABLE_s1_writedata                                        (mm_interconnect_0_spill_enable_s1_writedata),  //                                                           .writedata
		.SPILL_ENABLE_s1_chipselect                                       (mm_interconnect_0_spill_enable_s1_chipselect), //                                                           .chipselect
		.TICK_IN_s1_address                                               (mm_interconnect_0_tick_in_s1_address),         //                                                 TICK_IN_s1.address
		.TICK_IN_s1_write                                                 (mm_interconnect_0_tick_in_s1_write),           //                                                           .write
		.TICK_IN_s1_readdata                                              (mm_interconnect_0_tick_in_s1_readdata),        //                                                           .readdata
		.TICK_IN_s1_writedata                                             (mm_interconnect_0_tick_in_s1_writedata),       //                                                           .writedata
		.TICK_IN_s1_chipselect                                            (mm_interconnect_0_tick_in_s1_chipselect),      //                                                           .chipselect
		.TICK_OUT_s1_address                                              (mm_interconnect_0_tick_out_s1_address),        //                                                TICK_OUT_s1.address
		.TICK_OUT_s1_readdata                                             (mm_interconnect_0_tick_out_s1_readdata),       //                                                           .readdata
		.TIME_IN_s1_address                                               (mm_interconnect_0_time_in_s1_address),         //                                                 TIME_IN_s1.address
		.TIME_IN_s1_write                                                 (mm_interconnect_0_time_in_s1_write),           //                                                           .write
		.TIME_IN_s1_readdata                                              (mm_interconnect_0_time_in_s1_readdata),        //                                                           .readdata
		.TIME_IN_s1_writedata                                             (mm_interconnect_0_time_in_s1_writedata),       //                                                           .writedata
		.TIME_IN_s1_chipselect                                            (mm_interconnect_0_time_in_s1_chipselect),      //                                                           .chipselect
		.TIME_OUT_s1_address                                              (mm_interconnect_0_time_out_s1_address),        //                                                TIME_OUT_s1.address
		.TIME_OUT_s1_readdata                                             (mm_interconnect_0_time_out_s1_readdata),       //                                                           .readdata
		.TX_CLK_DIV_s1_address                                            (mm_interconnect_0_tx_clk_div_s1_address),      //                                              TX_CLK_DIV_s1.address
		.TX_CLK_DIV_s1_write                                              (mm_interconnect_0_tx_clk_div_s1_write),        //                                                           .write
		.TX_CLK_DIV_s1_readdata                                           (mm_interconnect_0_tx_clk_div_s1_readdata),     //                                                           .readdata
		.TX_CLK_DIV_s1_writedata                                          (mm_interconnect_0_tx_clk_div_s1_writedata),    //                                                           .writedata
		.TX_CLK_DIV_s1_chipselect                                         (mm_interconnect_0_tx_clk_div_s1_chipselect),   //                                                           .chipselect
		.TX_FULL_s1_address                                               (mm_interconnect_0_tx_full_s1_address),         //                                                 TX_FULL_s1.address
		.TX_FULL_s1_readdata                                              (mm_interconnect_0_tx_full_s1_readdata),        //                                                           .readdata
		.WR_DATA_s1_address                                               (mm_interconnect_0_wr_data_s1_address),         //                                                 WR_DATA_s1.address
		.WR_DATA_s1_write                                                 (mm_interconnect_0_wr_data_s1_write),           //                                                           .write
		.WR_DATA_s1_readdata                                              (mm_interconnect_0_wr_data_s1_readdata),        //                                                           .readdata
		.WR_DATA_s1_writedata                                             (mm_interconnect_0_wr_data_s1_writedata),       //                                                           .writedata
		.WR_DATA_s1_chipselect                                            (mm_interconnect_0_wr_data_s1_chipselect)       //                                                           .chipselect
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~hps_0_h2f_reset_reset),             // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
