// ulight_fifo.v

// Generated using ACDS version 17.1 593

`timescale 1 ps / 1 ps
module ulight_fifo (
		output wire        auto_start_external_connection_export,           //           auto_start_external_connection.export
		input  wire        clk_clk,                                         //                                      clk.clk
		output wire [2:0]  clock_sel_external_connection_export,            //            clock_sel_external_connection.export
		input  wire [5:0]  counter_rx_fifo_external_connection_export,      //      counter_rx_fifo_external_connection.export
		input  wire [5:0]  counter_tx_fifo_external_connection_export,      //      counter_tx_fifo_external_connection.export
		input  wire [8:0]  data_flag_rx_external_connection_export,         //         data_flag_rx_external_connection.export
		input  wire [13:0] data_info_external_connection_export,            //            data_info_external_connection.export
		output wire        data_read_en_rx_external_connection_export,      //      data_read_en_rx_external_connection.export
		input  wire        fifo_empty_rx_status_external_connection_export, // fifo_empty_rx_status_external_connection.export
		input  wire        fifo_empty_tx_status_external_connection_export, // fifo_empty_tx_status_external_connection.export
		input  wire        fifo_full_rx_status_external_connection_export,  //  fifo_full_rx_status_external_connection.export
		input  wire        fifo_full_tx_status_external_connection_export,  //  fifo_full_tx_status_external_connection.export
		input  wire [5:0]  fsm_info_external_connection_export,             //             fsm_info_external_connection.export
		output wire [4:0]  led_pio_test_external_connection_export,         //         led_pio_test_external_connection.export
		output wire        link_disable_external_connection_export,         //         link_disable_external_connection.export
		output wire        link_start_external_connection_export,           //           link_start_external_connection.export
		output wire [12:0] memory_mem_a,                                    //                                   memory.mem_a
		output wire [2:0]  memory_mem_ba,                                   //                                         .mem_ba
		output wire        memory_mem_ck,                                   //                                         .mem_ck
		output wire        memory_mem_ck_n,                                 //                                         .mem_ck_n
		output wire        memory_mem_cke,                                  //                                         .mem_cke
		output wire        memory_mem_cs_n,                                 //                                         .mem_cs_n
		output wire        memory_mem_ras_n,                                //                                         .mem_ras_n
		output wire        memory_mem_cas_n,                                //                                         .mem_cas_n
		output wire        memory_mem_we_n,                                 //                                         .mem_we_n
		output wire        memory_mem_reset_n,                              //                                         .mem_reset_n
		inout  wire [7:0]  memory_mem_dq,                                   //                                         .mem_dq
		inout  wire        memory_mem_dqs,                                  //                                         .mem_dqs
		inout  wire        memory_mem_dqs_n,                                //                                         .mem_dqs_n
		output wire        memory_mem_odt,                                  //                                         .mem_odt
		output wire        memory_mem_dm,                                   //                                         .mem_dm
		input  wire        memory_oct_rzqin,                                //                                         .oct_rzqin
		output wire        pll_0_locked_export,                             //                             pll_0_locked.export
		output wire        pll_0_outclk0_clk,                               //                            pll_0_outclk0.clk
		input  wire        reset_reset_n,                                   //                                    reset.reset_n
		input  wire        timecode_ready_rx_external_connection_export,    //    timecode_ready_rx_external_connection.export
		input  wire [7:0]  timecode_rx_external_connection_export,          //          timecode_rx_external_connection.export
		output wire [7:0]  timecode_tx_data_external_connection_export,     //     timecode_tx_data_external_connection.export
		output wire        timecode_tx_enable_external_connection_export,   //   timecode_tx_enable_external_connection.export
		input  wire        timecode_tx_ready_external_connection_export,    //    timecode_tx_ready_external_connection.export
		output wire [8:0]  write_data_fifo_tx_external_connection_export,   //   write_data_fifo_tx_external_connection.export
		output wire        write_en_tx_external_connection_export           //          write_en_tx_external_connection.export
	);

	wire   [1:0] hps_0_h2f_axi_master_awburst;                       // hps_0:h2f_AWBURST -> mm_interconnect_0:hps_0_h2f_axi_master_awburst
	wire   [3:0] hps_0_h2f_axi_master_arlen;                         // hps_0:h2f_ARLEN -> mm_interconnect_0:hps_0_h2f_axi_master_arlen
	wire   [3:0] hps_0_h2f_axi_master_wstrb;                         // hps_0:h2f_WSTRB -> mm_interconnect_0:hps_0_h2f_axi_master_wstrb
	wire         hps_0_h2f_axi_master_wready;                        // mm_interconnect_0:hps_0_h2f_axi_master_wready -> hps_0:h2f_WREADY
	wire  [11:0] hps_0_h2f_axi_master_rid;                           // mm_interconnect_0:hps_0_h2f_axi_master_rid -> hps_0:h2f_RID
	wire         hps_0_h2f_axi_master_rready;                        // hps_0:h2f_RREADY -> mm_interconnect_0:hps_0_h2f_axi_master_rready
	wire   [3:0] hps_0_h2f_axi_master_awlen;                         // hps_0:h2f_AWLEN -> mm_interconnect_0:hps_0_h2f_axi_master_awlen
	wire  [11:0] hps_0_h2f_axi_master_wid;                           // hps_0:h2f_WID -> mm_interconnect_0:hps_0_h2f_axi_master_wid
	wire   [3:0] hps_0_h2f_axi_master_arcache;                       // hps_0:h2f_ARCACHE -> mm_interconnect_0:hps_0_h2f_axi_master_arcache
	wire         hps_0_h2f_axi_master_wvalid;                        // hps_0:h2f_WVALID -> mm_interconnect_0:hps_0_h2f_axi_master_wvalid
	wire  [29:0] hps_0_h2f_axi_master_araddr;                        // hps_0:h2f_ARADDR -> mm_interconnect_0:hps_0_h2f_axi_master_araddr
	wire   [2:0] hps_0_h2f_axi_master_arprot;                        // hps_0:h2f_ARPROT -> mm_interconnect_0:hps_0_h2f_axi_master_arprot
	wire   [2:0] hps_0_h2f_axi_master_awprot;                        // hps_0:h2f_AWPROT -> mm_interconnect_0:hps_0_h2f_axi_master_awprot
	wire  [31:0] hps_0_h2f_axi_master_wdata;                         // hps_0:h2f_WDATA -> mm_interconnect_0:hps_0_h2f_axi_master_wdata
	wire         hps_0_h2f_axi_master_arvalid;                       // hps_0:h2f_ARVALID -> mm_interconnect_0:hps_0_h2f_axi_master_arvalid
	wire   [3:0] hps_0_h2f_axi_master_awcache;                       // hps_0:h2f_AWCACHE -> mm_interconnect_0:hps_0_h2f_axi_master_awcache
	wire  [11:0] hps_0_h2f_axi_master_arid;                          // hps_0:h2f_ARID -> mm_interconnect_0:hps_0_h2f_axi_master_arid
	wire   [1:0] hps_0_h2f_axi_master_arlock;                        // hps_0:h2f_ARLOCK -> mm_interconnect_0:hps_0_h2f_axi_master_arlock
	wire   [1:0] hps_0_h2f_axi_master_awlock;                        // hps_0:h2f_AWLOCK -> mm_interconnect_0:hps_0_h2f_axi_master_awlock
	wire  [29:0] hps_0_h2f_axi_master_awaddr;                        // hps_0:h2f_AWADDR -> mm_interconnect_0:hps_0_h2f_axi_master_awaddr
	wire   [1:0] hps_0_h2f_axi_master_bresp;                         // mm_interconnect_0:hps_0_h2f_axi_master_bresp -> hps_0:h2f_BRESP
	wire         hps_0_h2f_axi_master_arready;                       // mm_interconnect_0:hps_0_h2f_axi_master_arready -> hps_0:h2f_ARREADY
	wire  [31:0] hps_0_h2f_axi_master_rdata;                         // mm_interconnect_0:hps_0_h2f_axi_master_rdata -> hps_0:h2f_RDATA
	wire         hps_0_h2f_axi_master_awready;                       // mm_interconnect_0:hps_0_h2f_axi_master_awready -> hps_0:h2f_AWREADY
	wire   [1:0] hps_0_h2f_axi_master_arburst;                       // hps_0:h2f_ARBURST -> mm_interconnect_0:hps_0_h2f_axi_master_arburst
	wire   [2:0] hps_0_h2f_axi_master_arsize;                        // hps_0:h2f_ARSIZE -> mm_interconnect_0:hps_0_h2f_axi_master_arsize
	wire         hps_0_h2f_axi_master_bready;                        // hps_0:h2f_BREADY -> mm_interconnect_0:hps_0_h2f_axi_master_bready
	wire         hps_0_h2f_axi_master_rlast;                         // mm_interconnect_0:hps_0_h2f_axi_master_rlast -> hps_0:h2f_RLAST
	wire         hps_0_h2f_axi_master_wlast;                         // hps_0:h2f_WLAST -> mm_interconnect_0:hps_0_h2f_axi_master_wlast
	wire   [1:0] hps_0_h2f_axi_master_rresp;                         // mm_interconnect_0:hps_0_h2f_axi_master_rresp -> hps_0:h2f_RRESP
	wire  [11:0] hps_0_h2f_axi_master_awid;                          // hps_0:h2f_AWID -> mm_interconnect_0:hps_0_h2f_axi_master_awid
	wire  [11:0] hps_0_h2f_axi_master_bid;                           // mm_interconnect_0:hps_0_h2f_axi_master_bid -> hps_0:h2f_BID
	wire         hps_0_h2f_axi_master_bvalid;                        // mm_interconnect_0:hps_0_h2f_axi_master_bvalid -> hps_0:h2f_BVALID
	wire   [2:0] hps_0_h2f_axi_master_awsize;                        // hps_0:h2f_AWSIZE -> mm_interconnect_0:hps_0_h2f_axi_master_awsize
	wire         hps_0_h2f_axi_master_awvalid;                       // hps_0:h2f_AWVALID -> mm_interconnect_0:hps_0_h2f_axi_master_awvalid
	wire         hps_0_h2f_axi_master_rvalid;                        // mm_interconnect_0:hps_0_h2f_axi_master_rvalid -> hps_0:h2f_RVALID
	wire         mm_interconnect_0_led_pio_test_s1_chipselect;       // mm_interconnect_0:led_pio_test_s1_chipselect -> led_pio_test:chipselect
	wire  [31:0] mm_interconnect_0_led_pio_test_s1_readdata;         // led_pio_test:readdata -> mm_interconnect_0:led_pio_test_s1_readdata
	wire   [1:0] mm_interconnect_0_led_pio_test_s1_address;          // mm_interconnect_0:led_pio_test_s1_address -> led_pio_test:address
	wire         mm_interconnect_0_led_pio_test_s1_write;            // mm_interconnect_0:led_pio_test_s1_write -> led_pio_test:write_n
	wire  [31:0] mm_interconnect_0_led_pio_test_s1_writedata;        // mm_interconnect_0:led_pio_test_s1_writedata -> led_pio_test:writedata
	wire  [31:0] mm_interconnect_0_timecode_rx_s1_readdata;          // timecode_rx:readdata -> mm_interconnect_0:timecode_rx_s1_readdata
	wire   [1:0] mm_interconnect_0_timecode_rx_s1_address;           // mm_interconnect_0:timecode_rx_s1_address -> timecode_rx:address
	wire  [31:0] mm_interconnect_0_timecode_ready_rx_s1_readdata;    // timecode_ready_rx:readdata -> mm_interconnect_0:timecode_ready_rx_s1_readdata
	wire   [1:0] mm_interconnect_0_timecode_ready_rx_s1_address;     // mm_interconnect_0:timecode_ready_rx_s1_address -> timecode_ready_rx:address
	wire  [31:0] mm_interconnect_0_data_flag_rx_s1_readdata;         // data_flag_rx:readdata -> mm_interconnect_0:data_flag_rx_s1_readdata
	wire   [1:0] mm_interconnect_0_data_flag_rx_s1_address;          // mm_interconnect_0:data_flag_rx_s1_address -> data_flag_rx:address
	wire         mm_interconnect_0_data_read_en_rx_s1_chipselect;    // mm_interconnect_0:data_read_en_rx_s1_chipselect -> data_read_en_rx:chipselect
	wire  [31:0] mm_interconnect_0_data_read_en_rx_s1_readdata;      // data_read_en_rx:readdata -> mm_interconnect_0:data_read_en_rx_s1_readdata
	wire   [1:0] mm_interconnect_0_data_read_en_rx_s1_address;       // mm_interconnect_0:data_read_en_rx_s1_address -> data_read_en_rx:address
	wire         mm_interconnect_0_data_read_en_rx_s1_write;         // mm_interconnect_0:data_read_en_rx_s1_write -> data_read_en_rx:write_n
	wire  [31:0] mm_interconnect_0_data_read_en_rx_s1_writedata;     // mm_interconnect_0:data_read_en_rx_s1_writedata -> data_read_en_rx:writedata
	wire  [31:0] mm_interconnect_0_fifo_full_rx_status_s1_readdata;  // fifo_full_rx_status:readdata -> mm_interconnect_0:fifo_full_rx_status_s1_readdata
	wire   [1:0] mm_interconnect_0_fifo_full_rx_status_s1_address;   // mm_interconnect_0:fifo_full_rx_status_s1_address -> fifo_full_rx_status:address
	wire  [31:0] mm_interconnect_0_fifo_empty_rx_status_s1_readdata; // fifo_empty_rx_status:readdata -> mm_interconnect_0:fifo_empty_rx_status_s1_readdata
	wire   [1:0] mm_interconnect_0_fifo_empty_rx_status_s1_address;  // mm_interconnect_0:fifo_empty_rx_status_s1_address -> fifo_empty_rx_status:address
	wire         mm_interconnect_0_link_start_s1_chipselect;         // mm_interconnect_0:link_start_s1_chipselect -> link_start:chipselect
	wire  [31:0] mm_interconnect_0_link_start_s1_readdata;           // link_start:readdata -> mm_interconnect_0:link_start_s1_readdata
	wire   [1:0] mm_interconnect_0_link_start_s1_address;            // mm_interconnect_0:link_start_s1_address -> link_start:address
	wire         mm_interconnect_0_link_start_s1_write;              // mm_interconnect_0:link_start_s1_write -> link_start:write_n
	wire  [31:0] mm_interconnect_0_link_start_s1_writedata;          // mm_interconnect_0:link_start_s1_writedata -> link_start:writedata
	wire         mm_interconnect_0_auto_start_s1_chipselect;         // mm_interconnect_0:auto_start_s1_chipselect -> auto_start:chipselect
	wire  [31:0] mm_interconnect_0_auto_start_s1_readdata;           // auto_start:readdata -> mm_interconnect_0:auto_start_s1_readdata
	wire   [1:0] mm_interconnect_0_auto_start_s1_address;            // mm_interconnect_0:auto_start_s1_address -> auto_start:address
	wire         mm_interconnect_0_auto_start_s1_write;              // mm_interconnect_0:auto_start_s1_write -> auto_start:write_n
	wire  [31:0] mm_interconnect_0_auto_start_s1_writedata;          // mm_interconnect_0:auto_start_s1_writedata -> auto_start:writedata
	wire         mm_interconnect_0_link_disable_s1_chipselect;       // mm_interconnect_0:link_disable_s1_chipselect -> link_disable:chipselect
	wire  [31:0] mm_interconnect_0_link_disable_s1_readdata;         // link_disable:readdata -> mm_interconnect_0:link_disable_s1_readdata
	wire   [1:0] mm_interconnect_0_link_disable_s1_address;          // mm_interconnect_0:link_disable_s1_address -> link_disable:address
	wire         mm_interconnect_0_link_disable_s1_write;            // mm_interconnect_0:link_disable_s1_write -> link_disable:write_n
	wire  [31:0] mm_interconnect_0_link_disable_s1_writedata;        // mm_interconnect_0:link_disable_s1_writedata -> link_disable:writedata
	wire         mm_interconnect_0_write_data_fifo_tx_s1_chipselect; // mm_interconnect_0:write_data_fifo_tx_s1_chipselect -> write_data_fifo_tx:chipselect
	wire  [31:0] mm_interconnect_0_write_data_fifo_tx_s1_readdata;   // write_data_fifo_tx:readdata -> mm_interconnect_0:write_data_fifo_tx_s1_readdata
	wire   [1:0] mm_interconnect_0_write_data_fifo_tx_s1_address;    // mm_interconnect_0:write_data_fifo_tx_s1_address -> write_data_fifo_tx:address
	wire         mm_interconnect_0_write_data_fifo_tx_s1_write;      // mm_interconnect_0:write_data_fifo_tx_s1_write -> write_data_fifo_tx:write_n
	wire  [31:0] mm_interconnect_0_write_data_fifo_tx_s1_writedata;  // mm_interconnect_0:write_data_fifo_tx_s1_writedata -> write_data_fifo_tx:writedata
	wire         mm_interconnect_0_write_en_tx_s1_chipselect;        // mm_interconnect_0:write_en_tx_s1_chipselect -> write_en_tx:chipselect
	wire  [31:0] mm_interconnect_0_write_en_tx_s1_readdata;          // write_en_tx:readdata -> mm_interconnect_0:write_en_tx_s1_readdata
	wire   [1:0] mm_interconnect_0_write_en_tx_s1_address;           // mm_interconnect_0:write_en_tx_s1_address -> write_en_tx:address
	wire         mm_interconnect_0_write_en_tx_s1_write;             // mm_interconnect_0:write_en_tx_s1_write -> write_en_tx:write_n
	wire  [31:0] mm_interconnect_0_write_en_tx_s1_writedata;         // mm_interconnect_0:write_en_tx_s1_writedata -> write_en_tx:writedata
	wire  [31:0] mm_interconnect_0_fifo_full_tx_status_s1_readdata;  // fifo_full_tx_status:readdata -> mm_interconnect_0:fifo_full_tx_status_s1_readdata
	wire   [1:0] mm_interconnect_0_fifo_full_tx_status_s1_address;   // mm_interconnect_0:fifo_full_tx_status_s1_address -> fifo_full_tx_status:address
	wire  [31:0] mm_interconnect_0_fifo_empty_tx_status_s1_readdata; // fifo_empty_tx_status:readdata -> mm_interconnect_0:fifo_empty_tx_status_s1_readdata
	wire   [1:0] mm_interconnect_0_fifo_empty_tx_status_s1_address;  // mm_interconnect_0:fifo_empty_tx_status_s1_address -> fifo_empty_tx_status:address
	wire         mm_interconnect_0_timecode_tx_data_s1_chipselect;   // mm_interconnect_0:timecode_tx_data_s1_chipselect -> timecode_tx_data:chipselect
	wire  [31:0] mm_interconnect_0_timecode_tx_data_s1_readdata;     // timecode_tx_data:readdata -> mm_interconnect_0:timecode_tx_data_s1_readdata
	wire   [1:0] mm_interconnect_0_timecode_tx_data_s1_address;      // mm_interconnect_0:timecode_tx_data_s1_address -> timecode_tx_data:address
	wire         mm_interconnect_0_timecode_tx_data_s1_write;        // mm_interconnect_0:timecode_tx_data_s1_write -> timecode_tx_data:write_n
	wire  [31:0] mm_interconnect_0_timecode_tx_data_s1_writedata;    // mm_interconnect_0:timecode_tx_data_s1_writedata -> timecode_tx_data:writedata
	wire         mm_interconnect_0_timecode_tx_enable_s1_chipselect; // mm_interconnect_0:timecode_tx_enable_s1_chipselect -> timecode_tx_enable:chipselect
	wire  [31:0] mm_interconnect_0_timecode_tx_enable_s1_readdata;   // timecode_tx_enable:readdata -> mm_interconnect_0:timecode_tx_enable_s1_readdata
	wire   [1:0] mm_interconnect_0_timecode_tx_enable_s1_address;    // mm_interconnect_0:timecode_tx_enable_s1_address -> timecode_tx_enable:address
	wire         mm_interconnect_0_timecode_tx_enable_s1_write;      // mm_interconnect_0:timecode_tx_enable_s1_write -> timecode_tx_enable:write_n
	wire  [31:0] mm_interconnect_0_timecode_tx_enable_s1_writedata;  // mm_interconnect_0:timecode_tx_enable_s1_writedata -> timecode_tx_enable:writedata
	wire  [31:0] mm_interconnect_0_timecode_tx_ready_s1_readdata;    // timecode_tx_ready:readdata -> mm_interconnect_0:timecode_tx_ready_s1_readdata
	wire   [1:0] mm_interconnect_0_timecode_tx_ready_s1_address;     // mm_interconnect_0:timecode_tx_ready_s1_address -> timecode_tx_ready:address
	wire  [31:0] mm_interconnect_0_data_info_s1_readdata;            // data_info:readdata -> mm_interconnect_0:data_info_s1_readdata
	wire   [1:0] mm_interconnect_0_data_info_s1_address;             // mm_interconnect_0:data_info_s1_address -> data_info:address
	wire         mm_interconnect_0_clock_sel_s1_chipselect;          // mm_interconnect_0:clock_sel_s1_chipselect -> clock_sel:chipselect
	wire  [31:0] mm_interconnect_0_clock_sel_s1_readdata;            // clock_sel:readdata -> mm_interconnect_0:clock_sel_s1_readdata
	wire   [1:0] mm_interconnect_0_clock_sel_s1_address;             // mm_interconnect_0:clock_sel_s1_address -> clock_sel:address
	wire         mm_interconnect_0_clock_sel_s1_write;               // mm_interconnect_0:clock_sel_s1_write -> clock_sel:write_n
	wire  [31:0] mm_interconnect_0_clock_sel_s1_writedata;           // mm_interconnect_0:clock_sel_s1_writedata -> clock_sel:writedata
	wire  [31:0] mm_interconnect_0_fsm_info_s1_readdata;             // fsm_info:readdata -> mm_interconnect_0:fsm_info_s1_readdata
	wire   [1:0] mm_interconnect_0_fsm_info_s1_address;              // mm_interconnect_0:fsm_info_s1_address -> fsm_info:address
	wire  [31:0] mm_interconnect_0_counter_tx_fifo_s1_readdata;      // counter_tx_fifo:readdata -> mm_interconnect_0:counter_tx_fifo_s1_readdata
	wire   [1:0] mm_interconnect_0_counter_tx_fifo_s1_address;       // mm_interconnect_0:counter_tx_fifo_s1_address -> counter_tx_fifo:address
	wire  [31:0] mm_interconnect_0_counter_rx_fifo_s1_readdata;      // counter_rx_fifo:readdata -> mm_interconnect_0:counter_rx_fifo_s1_readdata
	wire   [1:0] mm_interconnect_0_counter_rx_fifo_s1_address;       // mm_interconnect_0:counter_rx_fifo_s1_address -> counter_rx_fifo:address
	wire         rst_controller_reset_out_reset;                     // rst_controller:reset_out -> [auto_start:reset_n, clock_sel:reset_n, counter_rx_fifo:reset_n, counter_tx_fifo:reset_n, data_flag_rx:reset_n, data_info:reset_n, data_read_en_rx:reset_n, fifo_empty_rx_status:reset_n, fifo_empty_tx_status:reset_n, fifo_full_rx_status:reset_n, fifo_full_tx_status:reset_n, fsm_info:reset_n, led_pio_test:reset_n, link_disable:reset_n, link_start:reset_n, mm_interconnect_0:led_pio_test_reset_reset_bridge_in_reset_reset, timecode_ready_rx:reset_n, timecode_rx:reset_n, timecode_tx_data:reset_n, timecode_tx_enable:reset_n, timecode_tx_ready:reset_n, write_data_fifo_tx:reset_n, write_en_tx:reset_n]
	wire         rst_controller_001_reset_out_reset;                 // rst_controller_001:reset_out -> mm_interconnect_0:hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset
	wire         hps_0_h2f_reset_reset;                              // hps_0:h2f_rst_n -> rst_controller_001:reset_in0

	ulight_fifo_auto_start auto_start (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_auto_start_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_auto_start_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_auto_start_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_auto_start_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_auto_start_s1_readdata),   //                    .readdata
		.out_port   (auto_start_external_connection_export)       // external_connection.export
	);

	ulight_fifo_clock_sel clock_sel (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_clock_sel_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_clock_sel_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_clock_sel_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_clock_sel_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_clock_sel_s1_readdata),   //                    .readdata
		.out_port   (clock_sel_external_connection_export)       // external_connection.export
	);

	ulight_fifo_counter_rx_fifo counter_rx_fifo (
		.clk      (clk_clk),                                       //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address  (mm_interconnect_0_counter_rx_fifo_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_counter_rx_fifo_s1_readdata), //                    .readdata
		.in_port  (counter_rx_fifo_external_connection_export)     // external_connection.export
	);

	ulight_fifo_counter_rx_fifo counter_tx_fifo (
		.clk      (clk_clk),                                       //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address  (mm_interconnect_0_counter_tx_fifo_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_counter_tx_fifo_s1_readdata), //                    .readdata
		.in_port  (counter_tx_fifo_external_connection_export)     // external_connection.export
	);

	ulight_fifo_data_flag_rx data_flag_rx (
		.clk      (clk_clk),                                    //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_0_data_flag_rx_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_data_flag_rx_s1_readdata), //                    .readdata
		.in_port  (data_flag_rx_external_connection_export)     // external_connection.export
	);

	ulight_fifo_data_info data_info (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address  (mm_interconnect_0_data_info_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_data_info_s1_readdata), //                    .readdata
		.in_port  (data_info_external_connection_export)     // external_connection.export
	);

	ulight_fifo_auto_start data_read_en_rx (
		.clk        (clk_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_data_read_en_rx_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_data_read_en_rx_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_data_read_en_rx_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_data_read_en_rx_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_data_read_en_rx_s1_readdata),   //                    .readdata
		.out_port   (data_read_en_rx_external_connection_export)       // external_connection.export
	);

	ulight_fifo_fifo_empty_rx_status fifo_empty_rx_status (
		.clk      (clk_clk),                                            //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                    //               reset.reset_n
		.address  (mm_interconnect_0_fifo_empty_rx_status_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_fifo_empty_rx_status_s1_readdata), //                    .readdata
		.in_port  (fifo_empty_rx_status_external_connection_export)     // external_connection.export
	);

	ulight_fifo_fifo_empty_rx_status fifo_empty_tx_status (
		.clk      (clk_clk),                                            //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                    //               reset.reset_n
		.address  (mm_interconnect_0_fifo_empty_tx_status_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_fifo_empty_tx_status_s1_readdata), //                    .readdata
		.in_port  (fifo_empty_tx_status_external_connection_export)     // external_connection.export
	);

	ulight_fifo_fifo_empty_rx_status fifo_full_rx_status (
		.clk      (clk_clk),                                           //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address  (mm_interconnect_0_fifo_full_rx_status_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_fifo_full_rx_status_s1_readdata), //                    .readdata
		.in_port  (fifo_full_rx_status_external_connection_export)     // external_connection.export
	);

	ulight_fifo_fifo_empty_rx_status fifo_full_tx_status (
		.clk      (clk_clk),                                           //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address  (mm_interconnect_0_fifo_full_tx_status_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_fifo_full_tx_status_s1_readdata), //                    .readdata
		.in_port  (fifo_full_tx_status_external_connection_export)     // external_connection.export
	);

	ulight_fifo_counter_rx_fifo fsm_info (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_fsm_info_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_fsm_info_s1_readdata), //                    .readdata
		.in_port  (fsm_info_external_connection_export)     // external_connection.export
	);

	ulight_fifo_hps_0 #(
		.F2S_Width (0),
		.S2F_Width (1)
	) hps_0 (
		.mem_a       (memory_mem_a),                 //         memory.mem_a
		.mem_ba      (memory_mem_ba),                //               .mem_ba
		.mem_ck      (memory_mem_ck),                //               .mem_ck
		.mem_ck_n    (memory_mem_ck_n),              //               .mem_ck_n
		.mem_cke     (memory_mem_cke),               //               .mem_cke
		.mem_cs_n    (memory_mem_cs_n),              //               .mem_cs_n
		.mem_ras_n   (memory_mem_ras_n),             //               .mem_ras_n
		.mem_cas_n   (memory_mem_cas_n),             //               .mem_cas_n
		.mem_we_n    (memory_mem_we_n),              //               .mem_we_n
		.mem_reset_n (memory_mem_reset_n),           //               .mem_reset_n
		.mem_dq      (memory_mem_dq),                //               .mem_dq
		.mem_dqs     (memory_mem_dqs),               //               .mem_dqs
		.mem_dqs_n   (memory_mem_dqs_n),             //               .mem_dqs_n
		.mem_odt     (memory_mem_odt),               //               .mem_odt
		.mem_dm      (memory_mem_dm),                //               .mem_dm
		.oct_rzqin   (memory_oct_rzqin),             //               .oct_rzqin
		.h2f_rst_n   (hps_0_h2f_reset_reset),        //      h2f_reset.reset_n
		.h2f_axi_clk (clk_clk),                      //  h2f_axi_clock.clk
		.h2f_AWID    (hps_0_h2f_axi_master_awid),    // h2f_axi_master.awid
		.h2f_AWADDR  (hps_0_h2f_axi_master_awaddr),  //               .awaddr
		.h2f_AWLEN   (hps_0_h2f_axi_master_awlen),   //               .awlen
		.h2f_AWSIZE  (hps_0_h2f_axi_master_awsize),  //               .awsize
		.h2f_AWBURST (hps_0_h2f_axi_master_awburst), //               .awburst
		.h2f_AWLOCK  (hps_0_h2f_axi_master_awlock),  //               .awlock
		.h2f_AWCACHE (hps_0_h2f_axi_master_awcache), //               .awcache
		.h2f_AWPROT  (hps_0_h2f_axi_master_awprot),  //               .awprot
		.h2f_AWVALID (hps_0_h2f_axi_master_awvalid), //               .awvalid
		.h2f_AWREADY (hps_0_h2f_axi_master_awready), //               .awready
		.h2f_WID     (hps_0_h2f_axi_master_wid),     //               .wid
		.h2f_WDATA   (hps_0_h2f_axi_master_wdata),   //               .wdata
		.h2f_WSTRB   (hps_0_h2f_axi_master_wstrb),   //               .wstrb
		.h2f_WLAST   (hps_0_h2f_axi_master_wlast),   //               .wlast
		.h2f_WVALID  (hps_0_h2f_axi_master_wvalid),  //               .wvalid
		.h2f_WREADY  (hps_0_h2f_axi_master_wready),  //               .wready
		.h2f_BID     (hps_0_h2f_axi_master_bid),     //               .bid
		.h2f_BRESP   (hps_0_h2f_axi_master_bresp),   //               .bresp
		.h2f_BVALID  (hps_0_h2f_axi_master_bvalid),  //               .bvalid
		.h2f_BREADY  (hps_0_h2f_axi_master_bready),  //               .bready
		.h2f_ARID    (hps_0_h2f_axi_master_arid),    //               .arid
		.h2f_ARADDR  (hps_0_h2f_axi_master_araddr),  //               .araddr
		.h2f_ARLEN   (hps_0_h2f_axi_master_arlen),   //               .arlen
		.h2f_ARSIZE  (hps_0_h2f_axi_master_arsize),  //               .arsize
		.h2f_ARBURST (hps_0_h2f_axi_master_arburst), //               .arburst
		.h2f_ARLOCK  (hps_0_h2f_axi_master_arlock),  //               .arlock
		.h2f_ARCACHE (hps_0_h2f_axi_master_arcache), //               .arcache
		.h2f_ARPROT  (hps_0_h2f_axi_master_arprot),  //               .arprot
		.h2f_ARVALID (hps_0_h2f_axi_master_arvalid), //               .arvalid
		.h2f_ARREADY (hps_0_h2f_axi_master_arready), //               .arready
		.h2f_RID     (hps_0_h2f_axi_master_rid),     //               .rid
		.h2f_RDATA   (hps_0_h2f_axi_master_rdata),   //               .rdata
		.h2f_RRESP   (hps_0_h2f_axi_master_rresp),   //               .rresp
		.h2f_RLAST   (hps_0_h2f_axi_master_rlast),   //               .rlast
		.h2f_RVALID  (hps_0_h2f_axi_master_rvalid),  //               .rvalid
		.h2f_RREADY  (hps_0_h2f_axi_master_rready)   //               .rready
	);

	ulight_fifo_led_pio_test led_pio_test (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_led_pio_test_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_pio_test_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_pio_test_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_pio_test_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_pio_test_s1_readdata),   //                    .readdata
		.out_port   (led_pio_test_external_connection_export)       // external_connection.export
	);

	ulight_fifo_auto_start link_disable (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_link_disable_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_link_disable_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_link_disable_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_link_disable_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_link_disable_s1_readdata),   //                    .readdata
		.out_port   (link_disable_external_connection_export)       // external_connection.export
	);

	ulight_fifo_auto_start link_start (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_link_start_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_link_start_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_link_start_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_link_start_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_link_start_s1_readdata),   //                    .readdata
		.out_port   (link_start_external_connection_export)       // external_connection.export
	);

	ulight_fifo_pll_0 pll_0 (
		.refclk   (clk_clk),             //  refclk.clk
		.rst      (~reset_reset_n),      //   reset.reset
		.outclk_0 (pll_0_outclk0_clk),   // outclk0.clk
		.locked   (pll_0_locked_export), //  locked.export
		.refclk1  ()                     // refclk1.refclk1
	);

	ulight_fifo_fifo_empty_rx_status timecode_ready_rx (
		.clk      (clk_clk),                                         //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address  (mm_interconnect_0_timecode_ready_rx_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_timecode_ready_rx_s1_readdata), //                    .readdata
		.in_port  (timecode_ready_rx_external_connection_export)     // external_connection.export
	);

	ulight_fifo_timecode_rx timecode_rx (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_0_timecode_rx_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_timecode_rx_s1_readdata), //                    .readdata
		.in_port  (timecode_rx_external_connection_export)     // external_connection.export
	);

	ulight_fifo_timecode_tx_data timecode_tx_data (
		.clk        (clk_clk),                                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (mm_interconnect_0_timecode_tx_data_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_timecode_tx_data_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_timecode_tx_data_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_timecode_tx_data_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_timecode_tx_data_s1_readdata),   //                    .readdata
		.out_port   (timecode_tx_data_external_connection_export)       // external_connection.export
	);

	ulight_fifo_auto_start timecode_tx_enable (
		.clk        (clk_clk),                                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                    //               reset.reset_n
		.address    (mm_interconnect_0_timecode_tx_enable_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_timecode_tx_enable_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_timecode_tx_enable_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_timecode_tx_enable_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_timecode_tx_enable_s1_readdata),   //                    .readdata
		.out_port   (timecode_tx_enable_external_connection_export)       // external_connection.export
	);

	ulight_fifo_fifo_empty_rx_status timecode_tx_ready (
		.clk      (clk_clk),                                         //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address  (mm_interconnect_0_timecode_tx_ready_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_timecode_tx_ready_s1_readdata), //                    .readdata
		.in_port  (timecode_tx_ready_external_connection_export)     // external_connection.export
	);

	ulight_fifo_write_data_fifo_tx write_data_fifo_tx (
		.clk        (clk_clk),                                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                    //               reset.reset_n
		.address    (mm_interconnect_0_write_data_fifo_tx_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_write_data_fifo_tx_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_write_data_fifo_tx_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_write_data_fifo_tx_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_write_data_fifo_tx_s1_readdata),   //                    .readdata
		.out_port   (write_data_fifo_tx_external_connection_export)       // external_connection.export
	);

	ulight_fifo_auto_start write_en_tx (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_write_en_tx_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_write_en_tx_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_write_en_tx_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_write_en_tx_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_write_en_tx_s1_readdata),   //                    .readdata
		.out_port   (write_en_tx_external_connection_export)       // external_connection.export
	);

	ulight_fifo_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_h2f_axi_master_awid                                        (hps_0_h2f_axi_master_awid),                          //                                       hps_0_h2f_axi_master.awid
		.hps_0_h2f_axi_master_awaddr                                      (hps_0_h2f_axi_master_awaddr),                        //                                                           .awaddr
		.hps_0_h2f_axi_master_awlen                                       (hps_0_h2f_axi_master_awlen),                         //                                                           .awlen
		.hps_0_h2f_axi_master_awsize                                      (hps_0_h2f_axi_master_awsize),                        //                                                           .awsize
		.hps_0_h2f_axi_master_awburst                                     (hps_0_h2f_axi_master_awburst),                       //                                                           .awburst
		.hps_0_h2f_axi_master_awlock                                      (hps_0_h2f_axi_master_awlock),                        //                                                           .awlock
		.hps_0_h2f_axi_master_awcache                                     (hps_0_h2f_axi_master_awcache),                       //                                                           .awcache
		.hps_0_h2f_axi_master_awprot                                      (hps_0_h2f_axi_master_awprot),                        //                                                           .awprot
		.hps_0_h2f_axi_master_awvalid                                     (hps_0_h2f_axi_master_awvalid),                       //                                                           .awvalid
		.hps_0_h2f_axi_master_awready                                     (hps_0_h2f_axi_master_awready),                       //                                                           .awready
		.hps_0_h2f_axi_master_wid                                         (hps_0_h2f_axi_master_wid),                           //                                                           .wid
		.hps_0_h2f_axi_master_wdata                                       (hps_0_h2f_axi_master_wdata),                         //                                                           .wdata
		.hps_0_h2f_axi_master_wstrb                                       (hps_0_h2f_axi_master_wstrb),                         //                                                           .wstrb
		.hps_0_h2f_axi_master_wlast                                       (hps_0_h2f_axi_master_wlast),                         //                                                           .wlast
		.hps_0_h2f_axi_master_wvalid                                      (hps_0_h2f_axi_master_wvalid),                        //                                                           .wvalid
		.hps_0_h2f_axi_master_wready                                      (hps_0_h2f_axi_master_wready),                        //                                                           .wready
		.hps_0_h2f_axi_master_bid                                         (hps_0_h2f_axi_master_bid),                           //                                                           .bid
		.hps_0_h2f_axi_master_bresp                                       (hps_0_h2f_axi_master_bresp),                         //                                                           .bresp
		.hps_0_h2f_axi_master_bvalid                                      (hps_0_h2f_axi_master_bvalid),                        //                                                           .bvalid
		.hps_0_h2f_axi_master_bready                                      (hps_0_h2f_axi_master_bready),                        //                                                           .bready
		.hps_0_h2f_axi_master_arid                                        (hps_0_h2f_axi_master_arid),                          //                                                           .arid
		.hps_0_h2f_axi_master_araddr                                      (hps_0_h2f_axi_master_araddr),                        //                                                           .araddr
		.hps_0_h2f_axi_master_arlen                                       (hps_0_h2f_axi_master_arlen),                         //                                                           .arlen
		.hps_0_h2f_axi_master_arsize                                      (hps_0_h2f_axi_master_arsize),                        //                                                           .arsize
		.hps_0_h2f_axi_master_arburst                                     (hps_0_h2f_axi_master_arburst),                       //                                                           .arburst
		.hps_0_h2f_axi_master_arlock                                      (hps_0_h2f_axi_master_arlock),                        //                                                           .arlock
		.hps_0_h2f_axi_master_arcache                                     (hps_0_h2f_axi_master_arcache),                       //                                                           .arcache
		.hps_0_h2f_axi_master_arprot                                      (hps_0_h2f_axi_master_arprot),                        //                                                           .arprot
		.hps_0_h2f_axi_master_arvalid                                     (hps_0_h2f_axi_master_arvalid),                       //                                                           .arvalid
		.hps_0_h2f_axi_master_arready                                     (hps_0_h2f_axi_master_arready),                       //                                                           .arready
		.hps_0_h2f_axi_master_rid                                         (hps_0_h2f_axi_master_rid),                           //                                                           .rid
		.hps_0_h2f_axi_master_rdata                                       (hps_0_h2f_axi_master_rdata),                         //                                                           .rdata
		.hps_0_h2f_axi_master_rresp                                       (hps_0_h2f_axi_master_rresp),                         //                                                           .rresp
		.hps_0_h2f_axi_master_rlast                                       (hps_0_h2f_axi_master_rlast),                         //                                                           .rlast
		.hps_0_h2f_axi_master_rvalid                                      (hps_0_h2f_axi_master_rvalid),                        //                                                           .rvalid
		.hps_0_h2f_axi_master_rready                                      (hps_0_h2f_axi_master_rready),                        //                                                           .rready
		.clk_0_clk_clk                                                    (clk_clk),                                            //                                                  clk_0_clk.clk
		.hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                 // hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.led_pio_test_reset_reset_bridge_in_reset_reset                   (rst_controller_reset_out_reset),                     //                   led_pio_test_reset_reset_bridge_in_reset.reset
		.auto_start_s1_address                                            (mm_interconnect_0_auto_start_s1_address),            //                                              auto_start_s1.address
		.auto_start_s1_write                                              (mm_interconnect_0_auto_start_s1_write),              //                                                           .write
		.auto_start_s1_readdata                                           (mm_interconnect_0_auto_start_s1_readdata),           //                                                           .readdata
		.auto_start_s1_writedata                                          (mm_interconnect_0_auto_start_s1_writedata),          //                                                           .writedata
		.auto_start_s1_chipselect                                         (mm_interconnect_0_auto_start_s1_chipselect),         //                                                           .chipselect
		.clock_sel_s1_address                                             (mm_interconnect_0_clock_sel_s1_address),             //                                               clock_sel_s1.address
		.clock_sel_s1_write                                               (mm_interconnect_0_clock_sel_s1_write),               //                                                           .write
		.clock_sel_s1_readdata                                            (mm_interconnect_0_clock_sel_s1_readdata),            //                                                           .readdata
		.clock_sel_s1_writedata                                           (mm_interconnect_0_clock_sel_s1_writedata),           //                                                           .writedata
		.clock_sel_s1_chipselect                                          (mm_interconnect_0_clock_sel_s1_chipselect),          //                                                           .chipselect
		.counter_rx_fifo_s1_address                                       (mm_interconnect_0_counter_rx_fifo_s1_address),       //                                         counter_rx_fifo_s1.address
		.counter_rx_fifo_s1_readdata                                      (mm_interconnect_0_counter_rx_fifo_s1_readdata),      //                                                           .readdata
		.counter_tx_fifo_s1_address                                       (mm_interconnect_0_counter_tx_fifo_s1_address),       //                                         counter_tx_fifo_s1.address
		.counter_tx_fifo_s1_readdata                                      (mm_interconnect_0_counter_tx_fifo_s1_readdata),      //                                                           .readdata
		.data_flag_rx_s1_address                                          (mm_interconnect_0_data_flag_rx_s1_address),          //                                            data_flag_rx_s1.address
		.data_flag_rx_s1_readdata                                         (mm_interconnect_0_data_flag_rx_s1_readdata),         //                                                           .readdata
		.data_info_s1_address                                             (mm_interconnect_0_data_info_s1_address),             //                                               data_info_s1.address
		.data_info_s1_readdata                                            (mm_interconnect_0_data_info_s1_readdata),            //                                                           .readdata
		.data_read_en_rx_s1_address                                       (mm_interconnect_0_data_read_en_rx_s1_address),       //                                         data_read_en_rx_s1.address
		.data_read_en_rx_s1_write                                         (mm_interconnect_0_data_read_en_rx_s1_write),         //                                                           .write
		.data_read_en_rx_s1_readdata                                      (mm_interconnect_0_data_read_en_rx_s1_readdata),      //                                                           .readdata
		.data_read_en_rx_s1_writedata                                     (mm_interconnect_0_data_read_en_rx_s1_writedata),     //                                                           .writedata
		.data_read_en_rx_s1_chipselect                                    (mm_interconnect_0_data_read_en_rx_s1_chipselect),    //                                                           .chipselect
		.fifo_empty_rx_status_s1_address                                  (mm_interconnect_0_fifo_empty_rx_status_s1_address),  //                                    fifo_empty_rx_status_s1.address
		.fifo_empty_rx_status_s1_readdata                                 (mm_interconnect_0_fifo_empty_rx_status_s1_readdata), //                                                           .readdata
		.fifo_empty_tx_status_s1_address                                  (mm_interconnect_0_fifo_empty_tx_status_s1_address),  //                                    fifo_empty_tx_status_s1.address
		.fifo_empty_tx_status_s1_readdata                                 (mm_interconnect_0_fifo_empty_tx_status_s1_readdata), //                                                           .readdata
		.fifo_full_rx_status_s1_address                                   (mm_interconnect_0_fifo_full_rx_status_s1_address),   //                                     fifo_full_rx_status_s1.address
		.fifo_full_rx_status_s1_readdata                                  (mm_interconnect_0_fifo_full_rx_status_s1_readdata),  //                                                           .readdata
		.fifo_full_tx_status_s1_address                                   (mm_interconnect_0_fifo_full_tx_status_s1_address),   //                                     fifo_full_tx_status_s1.address
		.fifo_full_tx_status_s1_readdata                                  (mm_interconnect_0_fifo_full_tx_status_s1_readdata),  //                                                           .readdata
		.fsm_info_s1_address                                              (mm_interconnect_0_fsm_info_s1_address),              //                                                fsm_info_s1.address
		.fsm_info_s1_readdata                                             (mm_interconnect_0_fsm_info_s1_readdata),             //                                                           .readdata
		.led_pio_test_s1_address                                          (mm_interconnect_0_led_pio_test_s1_address),          //                                            led_pio_test_s1.address
		.led_pio_test_s1_write                                            (mm_interconnect_0_led_pio_test_s1_write),            //                                                           .write
		.led_pio_test_s1_readdata                                         (mm_interconnect_0_led_pio_test_s1_readdata),         //                                                           .readdata
		.led_pio_test_s1_writedata                                        (mm_interconnect_0_led_pio_test_s1_writedata),        //                                                           .writedata
		.led_pio_test_s1_chipselect                                       (mm_interconnect_0_led_pio_test_s1_chipselect),       //                                                           .chipselect
		.link_disable_s1_address                                          (mm_interconnect_0_link_disable_s1_address),          //                                            link_disable_s1.address
		.link_disable_s1_write                                            (mm_interconnect_0_link_disable_s1_write),            //                                                           .write
		.link_disable_s1_readdata                                         (mm_interconnect_0_link_disable_s1_readdata),         //                                                           .readdata
		.link_disable_s1_writedata                                        (mm_interconnect_0_link_disable_s1_writedata),        //                                                           .writedata
		.link_disable_s1_chipselect                                       (mm_interconnect_0_link_disable_s1_chipselect),       //                                                           .chipselect
		.link_start_s1_address                                            (mm_interconnect_0_link_start_s1_address),            //                                              link_start_s1.address
		.link_start_s1_write                                              (mm_interconnect_0_link_start_s1_write),              //                                                           .write
		.link_start_s1_readdata                                           (mm_interconnect_0_link_start_s1_readdata),           //                                                           .readdata
		.link_start_s1_writedata                                          (mm_interconnect_0_link_start_s1_writedata),          //                                                           .writedata
		.link_start_s1_chipselect                                         (mm_interconnect_0_link_start_s1_chipselect),         //                                                           .chipselect
		.timecode_ready_rx_s1_address                                     (mm_interconnect_0_timecode_ready_rx_s1_address),     //                                       timecode_ready_rx_s1.address
		.timecode_ready_rx_s1_readdata                                    (mm_interconnect_0_timecode_ready_rx_s1_readdata),    //                                                           .readdata
		.timecode_rx_s1_address                                           (mm_interconnect_0_timecode_rx_s1_address),           //                                             timecode_rx_s1.address
		.timecode_rx_s1_readdata                                          (mm_interconnect_0_timecode_rx_s1_readdata),          //                                                           .readdata
		.timecode_tx_data_s1_address                                      (mm_interconnect_0_timecode_tx_data_s1_address),      //                                        timecode_tx_data_s1.address
		.timecode_tx_data_s1_write                                        (mm_interconnect_0_timecode_tx_data_s1_write),        //                                                           .write
		.timecode_tx_data_s1_readdata                                     (mm_interconnect_0_timecode_tx_data_s1_readdata),     //                                                           .readdata
		.timecode_tx_data_s1_writedata                                    (mm_interconnect_0_timecode_tx_data_s1_writedata),    //                                                           .writedata
		.timecode_tx_data_s1_chipselect                                   (mm_interconnect_0_timecode_tx_data_s1_chipselect),   //                                                           .chipselect
		.timecode_tx_enable_s1_address                                    (mm_interconnect_0_timecode_tx_enable_s1_address),    //                                      timecode_tx_enable_s1.address
		.timecode_tx_enable_s1_write                                      (mm_interconnect_0_timecode_tx_enable_s1_write),      //                                                           .write
		.timecode_tx_enable_s1_readdata                                   (mm_interconnect_0_timecode_tx_enable_s1_readdata),   //                                                           .readdata
		.timecode_tx_enable_s1_writedata                                  (mm_interconnect_0_timecode_tx_enable_s1_writedata),  //                                                           .writedata
		.timecode_tx_enable_s1_chipselect                                 (mm_interconnect_0_timecode_tx_enable_s1_chipselect), //                                                           .chipselect
		.timecode_tx_ready_s1_address                                     (mm_interconnect_0_timecode_tx_ready_s1_address),     //                                       timecode_tx_ready_s1.address
		.timecode_tx_ready_s1_readdata                                    (mm_interconnect_0_timecode_tx_ready_s1_readdata),    //                                                           .readdata
		.write_data_fifo_tx_s1_address                                    (mm_interconnect_0_write_data_fifo_tx_s1_address),    //                                      write_data_fifo_tx_s1.address
		.write_data_fifo_tx_s1_write                                      (mm_interconnect_0_write_data_fifo_tx_s1_write),      //                                                           .write
		.write_data_fifo_tx_s1_readdata                                   (mm_interconnect_0_write_data_fifo_tx_s1_readdata),   //                                                           .readdata
		.write_data_fifo_tx_s1_writedata                                  (mm_interconnect_0_write_data_fifo_tx_s1_writedata),  //                                                           .writedata
		.write_data_fifo_tx_s1_chipselect                                 (mm_interconnect_0_write_data_fifo_tx_s1_chipselect), //                                                           .chipselect
		.write_en_tx_s1_address                                           (mm_interconnect_0_write_en_tx_s1_address),           //                                             write_en_tx_s1.address
		.write_en_tx_s1_write                                             (mm_interconnect_0_write_en_tx_s1_write),             //                                                           .write
		.write_en_tx_s1_readdata                                          (mm_interconnect_0_write_en_tx_s1_readdata),          //                                                           .readdata
		.write_en_tx_s1_writedata                                         (mm_interconnect_0_write_en_tx_s1_writedata),         //                                                           .writedata
		.write_en_tx_s1_chipselect                                        (mm_interconnect_0_write_en_tx_s1_chipselect)         //                                                           .chipselect
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~hps_0_h2f_reset_reset),             // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
