// spw_ulight_nofifo.v

// Generated using ACDS version 16.1 203

`timescale 1 ps / 1 ps
module spw_ulight_nofifo (
		output wire        auto_start_0_external_connection_export,      //      auto_start_0_external_connection.export
		output wire        auto_start_external_connection_export,        //        auto_start_external_connection.export
		input  wire        clk_clk,                                      //                                   clk.clk
		output wire [2:0]  clock_sel_external_connection_export,         //         clock_sel_external_connection.export
		output wire        credit_error_rx_0_external_connection_export, // credit_error_rx_0_external_connection.export
		output wire        credit_error_rx_external_connection_export,   //   credit_error_rx_external_connection.export
		output wire        data_en_to_w_0_external_connection_export,    //    data_en_to_w_0_external_connection.export
		output wire        data_en_to_w_external_connection_export,      //      data_en_to_w_external_connection.export
		input  wire [8:0]  data_rx_r_0_external_connection_export,       //       data_rx_r_0_external_connection.export
		input  wire [8:0]  data_rx_r_external_connection_export,         //         data_rx_r_external_connection.export
		input  wire        data_rx_ready_0_external_connection_export,   //   data_rx_ready_0_external_connection.export
		input  wire        data_rx_ready_external_connection_export,     //     data_rx_ready_external_connection.export
		input  wire        data_tx_ready_0_external_connection_export,   //   data_tx_ready_0_external_connection.export
		input  wire        data_tx_ready_external_connection_export,     //     data_tx_ready_external_connection.export
		output wire [8:0]  data_tx_to_w_0_external_connection_export,    //    data_tx_to_w_0_external_connection.export
		output wire [8:0]  data_tx_to_w_external_connection_export,      //      data_tx_to_w_external_connection.export
		input  wire [5:0]  fsm_info_0_external_connection_export,        //        fsm_info_0_external_connection.export
		input  wire [5:0]  fsm_info_external_connection_export,          //          fsm_info_external_connection.export
		output wire [5:0]  led_fpga_external_connection_export,          //          led_fpga_external_connection.export
		output wire        link_disable_0_external_connection_export,    //    link_disable_0_external_connection.export
		output wire        link_disable_external_connection_export,      //      link_disable_external_connection.export
		output wire        link_start_0_external_connection_export,      //      link_start_0_external_connection.export
		output wire        link_start_external_connection_export,        //        link_start_external_connection.export
		input  wire [13:0] monitor_a_external_connection_export,         //         monitor_a_external_connection.export
		input  wire [13:0] monitor_b_external_connection_export,         //         monitor_b_external_connection.export
		output wire        pll_tx_locked_export,                         //                         pll_tx_locked.export
		output wire        pll_tx_outclk0_clk,                           //                        pll_tx_outclk0.clk
		output wire        pll_tx_outclk1_clk,                           //                        pll_tx_outclk1.clk
		output wire        pll_tx_outclk2_clk,                           //                        pll_tx_outclk2.clk
		output wire        pll_tx_outclk3_clk,                           //                        pll_tx_outclk3.clk
		output wire        pll_tx_outclk4_clk,                           //                        pll_tx_outclk4.clk
		input  wire        reset_reset_n,                                //                                 reset.reset_n
		output wire        send_fct_now_0_external_connection_export,    //    send_fct_now_0_external_connection.export
		output wire        send_fct_now_external_connection_export,      //      send_fct_now_external_connection.export
		output wire        timec_en_to_tx_0_external_connection_export,  //  timec_en_to_tx_0_external_connection.export
		output wire        timec_en_to_tx_external_connection_export,    //    timec_en_to_tx_external_connection.export
		input  wire [7:0]  timec_rx_r_0_external_connection_export,      //      timec_rx_r_0_external_connection.export
		input  wire [7:0]  timec_rx_r_external_connection_export,        //        timec_rx_r_external_connection.export
		input  wire        timec_rx_ready_0_external_connection_export,  //  timec_rx_ready_0_external_connection.export
		input  wire        timec_rx_ready_external_connection_export,    //    timec_rx_ready_external_connection.export
		input  wire        timec_tx_ready_0_external_connection_export,  //  timec_tx_ready_0_external_connection.export
		input  wire        timec_tx_ready_external_connection_export,    //    timec_tx_ready_external_connection.export
		output wire [7:0]  timec_tx_to_w_0_external_connection_export,   //   timec_tx_to_w_0_external_connection.export
		output wire [7:0]  timec_tx_to_w_external_connection_export      //     timec_tx_to_w_external_connection.export
	);

	wire   [1:0] hps_0_h2f_axi_master_awburst;                      // hps_0:h2f_AWBURST -> mm_interconnect_0:hps_0_h2f_axi_master_awburst
	wire   [3:0] hps_0_h2f_axi_master_arlen;                        // hps_0:h2f_ARLEN -> mm_interconnect_0:hps_0_h2f_axi_master_arlen
	wire   [3:0] hps_0_h2f_axi_master_wstrb;                        // hps_0:h2f_WSTRB -> mm_interconnect_0:hps_0_h2f_axi_master_wstrb
	wire         hps_0_h2f_axi_master_wready;                       // mm_interconnect_0:hps_0_h2f_axi_master_wready -> hps_0:h2f_WREADY
	wire  [11:0] hps_0_h2f_axi_master_rid;                          // mm_interconnect_0:hps_0_h2f_axi_master_rid -> hps_0:h2f_RID
	wire         hps_0_h2f_axi_master_rready;                       // hps_0:h2f_RREADY -> mm_interconnect_0:hps_0_h2f_axi_master_rready
	wire   [3:0] hps_0_h2f_axi_master_awlen;                        // hps_0:h2f_AWLEN -> mm_interconnect_0:hps_0_h2f_axi_master_awlen
	wire  [11:0] hps_0_h2f_axi_master_wid;                          // hps_0:h2f_WID -> mm_interconnect_0:hps_0_h2f_axi_master_wid
	wire   [3:0] hps_0_h2f_axi_master_arcache;                      // hps_0:h2f_ARCACHE -> mm_interconnect_0:hps_0_h2f_axi_master_arcache
	wire         hps_0_h2f_axi_master_wvalid;                       // hps_0:h2f_WVALID -> mm_interconnect_0:hps_0_h2f_axi_master_wvalid
	wire  [29:0] hps_0_h2f_axi_master_araddr;                       // hps_0:h2f_ARADDR -> mm_interconnect_0:hps_0_h2f_axi_master_araddr
	wire   [2:0] hps_0_h2f_axi_master_arprot;                       // hps_0:h2f_ARPROT -> mm_interconnect_0:hps_0_h2f_axi_master_arprot
	wire   [2:0] hps_0_h2f_axi_master_awprot;                       // hps_0:h2f_AWPROT -> mm_interconnect_0:hps_0_h2f_axi_master_awprot
	wire  [31:0] hps_0_h2f_axi_master_wdata;                        // hps_0:h2f_WDATA -> mm_interconnect_0:hps_0_h2f_axi_master_wdata
	wire         hps_0_h2f_axi_master_arvalid;                      // hps_0:h2f_ARVALID -> mm_interconnect_0:hps_0_h2f_axi_master_arvalid
	wire   [3:0] hps_0_h2f_axi_master_awcache;                      // hps_0:h2f_AWCACHE -> mm_interconnect_0:hps_0_h2f_axi_master_awcache
	wire  [11:0] hps_0_h2f_axi_master_arid;                         // hps_0:h2f_ARID -> mm_interconnect_0:hps_0_h2f_axi_master_arid
	wire   [1:0] hps_0_h2f_axi_master_arlock;                       // hps_0:h2f_ARLOCK -> mm_interconnect_0:hps_0_h2f_axi_master_arlock
	wire   [1:0] hps_0_h2f_axi_master_awlock;                       // hps_0:h2f_AWLOCK -> mm_interconnect_0:hps_0_h2f_axi_master_awlock
	wire  [29:0] hps_0_h2f_axi_master_awaddr;                       // hps_0:h2f_AWADDR -> mm_interconnect_0:hps_0_h2f_axi_master_awaddr
	wire   [1:0] hps_0_h2f_axi_master_bresp;                        // mm_interconnect_0:hps_0_h2f_axi_master_bresp -> hps_0:h2f_BRESP
	wire         hps_0_h2f_axi_master_arready;                      // mm_interconnect_0:hps_0_h2f_axi_master_arready -> hps_0:h2f_ARREADY
	wire  [31:0] hps_0_h2f_axi_master_rdata;                        // mm_interconnect_0:hps_0_h2f_axi_master_rdata -> hps_0:h2f_RDATA
	wire         hps_0_h2f_axi_master_awready;                      // mm_interconnect_0:hps_0_h2f_axi_master_awready -> hps_0:h2f_AWREADY
	wire   [1:0] hps_0_h2f_axi_master_arburst;                      // hps_0:h2f_ARBURST -> mm_interconnect_0:hps_0_h2f_axi_master_arburst
	wire   [2:0] hps_0_h2f_axi_master_arsize;                       // hps_0:h2f_ARSIZE -> mm_interconnect_0:hps_0_h2f_axi_master_arsize
	wire         hps_0_h2f_axi_master_bready;                       // hps_0:h2f_BREADY -> mm_interconnect_0:hps_0_h2f_axi_master_bready
	wire         hps_0_h2f_axi_master_rlast;                        // mm_interconnect_0:hps_0_h2f_axi_master_rlast -> hps_0:h2f_RLAST
	wire         hps_0_h2f_axi_master_wlast;                        // hps_0:h2f_WLAST -> mm_interconnect_0:hps_0_h2f_axi_master_wlast
	wire   [1:0] hps_0_h2f_axi_master_rresp;                        // mm_interconnect_0:hps_0_h2f_axi_master_rresp -> hps_0:h2f_RRESP
	wire  [11:0] hps_0_h2f_axi_master_awid;                         // hps_0:h2f_AWID -> mm_interconnect_0:hps_0_h2f_axi_master_awid
	wire  [11:0] hps_0_h2f_axi_master_bid;                          // mm_interconnect_0:hps_0_h2f_axi_master_bid -> hps_0:h2f_BID
	wire         hps_0_h2f_axi_master_bvalid;                       // mm_interconnect_0:hps_0_h2f_axi_master_bvalid -> hps_0:h2f_BVALID
	wire   [2:0] hps_0_h2f_axi_master_awsize;                       // hps_0:h2f_AWSIZE -> mm_interconnect_0:hps_0_h2f_axi_master_awsize
	wire         hps_0_h2f_axi_master_awvalid;                      // hps_0:h2f_AWVALID -> mm_interconnect_0:hps_0_h2f_axi_master_awvalid
	wire         hps_0_h2f_axi_master_rvalid;                       // mm_interconnect_0:hps_0_h2f_axi_master_rvalid -> hps_0:h2f_RVALID
	wire         mm_interconnect_0_led_fpga_s1_chipselect;          // mm_interconnect_0:led_fpga_s1_chipselect -> led_fpga:chipselect
	wire  [31:0] mm_interconnect_0_led_fpga_s1_readdata;            // led_fpga:readdata -> mm_interconnect_0:led_fpga_s1_readdata
	wire   [1:0] mm_interconnect_0_led_fpga_s1_address;             // mm_interconnect_0:led_fpga_s1_address -> led_fpga:address
	wire         mm_interconnect_0_led_fpga_s1_write;               // mm_interconnect_0:led_fpga_s1_write -> led_fpga:write_n
	wire  [31:0] mm_interconnect_0_led_fpga_s1_writedata;           // mm_interconnect_0:led_fpga_s1_writedata -> led_fpga:writedata
	wire  [31:0] mm_interconnect_0_monitor_a_s1_readdata;           // MONITOR_A:readdata -> mm_interconnect_0:MONITOR_A_s1_readdata
	wire   [1:0] mm_interconnect_0_monitor_a_s1_address;            // mm_interconnect_0:MONITOR_A_s1_address -> MONITOR_A:address
	wire  [31:0] mm_interconnect_0_monitor_b_s1_readdata;           // MONITOR_B:readdata -> mm_interconnect_0:MONITOR_B_s1_readdata
	wire   [1:0] mm_interconnect_0_monitor_b_s1_address;            // mm_interconnect_0:MONITOR_B_s1_address -> MONITOR_B:address
	wire         mm_interconnect_0_auto_start_s1_chipselect;        // mm_interconnect_0:auto_start_s1_chipselect -> auto_start:chipselect
	wire  [31:0] mm_interconnect_0_auto_start_s1_readdata;          // auto_start:readdata -> mm_interconnect_0:auto_start_s1_readdata
	wire   [1:0] mm_interconnect_0_auto_start_s1_address;           // mm_interconnect_0:auto_start_s1_address -> auto_start:address
	wire         mm_interconnect_0_auto_start_s1_write;             // mm_interconnect_0:auto_start_s1_write -> auto_start:write_n
	wire  [31:0] mm_interconnect_0_auto_start_s1_writedata;         // mm_interconnect_0:auto_start_s1_writedata -> auto_start:writedata
	wire         mm_interconnect_0_auto_start_0_s1_chipselect;      // mm_interconnect_0:auto_start_0_s1_chipselect -> auto_start_0:chipselect
	wire  [31:0] mm_interconnect_0_auto_start_0_s1_readdata;        // auto_start_0:readdata -> mm_interconnect_0:auto_start_0_s1_readdata
	wire   [1:0] mm_interconnect_0_auto_start_0_s1_address;         // mm_interconnect_0:auto_start_0_s1_address -> auto_start_0:address
	wire         mm_interconnect_0_auto_start_0_s1_write;           // mm_interconnect_0:auto_start_0_s1_write -> auto_start_0:write_n
	wire  [31:0] mm_interconnect_0_auto_start_0_s1_writedata;       // mm_interconnect_0:auto_start_0_s1_writedata -> auto_start_0:writedata
	wire         mm_interconnect_0_clock_sel_s1_chipselect;         // mm_interconnect_0:clock_sel_s1_chipselect -> clock_sel:chipselect
	wire  [31:0] mm_interconnect_0_clock_sel_s1_readdata;           // clock_sel:readdata -> mm_interconnect_0:clock_sel_s1_readdata
	wire   [1:0] mm_interconnect_0_clock_sel_s1_address;            // mm_interconnect_0:clock_sel_s1_address -> clock_sel:address
	wire         mm_interconnect_0_clock_sel_s1_write;              // mm_interconnect_0:clock_sel_s1_write -> clock_sel:write_n
	wire  [31:0] mm_interconnect_0_clock_sel_s1_writedata;          // mm_interconnect_0:clock_sel_s1_writedata -> clock_sel:writedata
	wire         mm_interconnect_0_credit_error_rx_s1_chipselect;   // mm_interconnect_0:credit_error_rx_s1_chipselect -> credit_error_rx:chipselect
	wire  [31:0] mm_interconnect_0_credit_error_rx_s1_readdata;     // credit_error_rx:readdata -> mm_interconnect_0:credit_error_rx_s1_readdata
	wire   [1:0] mm_interconnect_0_credit_error_rx_s1_address;      // mm_interconnect_0:credit_error_rx_s1_address -> credit_error_rx:address
	wire         mm_interconnect_0_credit_error_rx_s1_write;        // mm_interconnect_0:credit_error_rx_s1_write -> credit_error_rx:write_n
	wire  [31:0] mm_interconnect_0_credit_error_rx_s1_writedata;    // mm_interconnect_0:credit_error_rx_s1_writedata -> credit_error_rx:writedata
	wire         mm_interconnect_0_credit_error_rx_0_s1_chipselect; // mm_interconnect_0:credit_error_rx_0_s1_chipselect -> credit_error_rx_0:chipselect
	wire  [31:0] mm_interconnect_0_credit_error_rx_0_s1_readdata;   // credit_error_rx_0:readdata -> mm_interconnect_0:credit_error_rx_0_s1_readdata
	wire   [1:0] mm_interconnect_0_credit_error_rx_0_s1_address;    // mm_interconnect_0:credit_error_rx_0_s1_address -> credit_error_rx_0:address
	wire         mm_interconnect_0_credit_error_rx_0_s1_write;      // mm_interconnect_0:credit_error_rx_0_s1_write -> credit_error_rx_0:write_n
	wire  [31:0] mm_interconnect_0_credit_error_rx_0_s1_writedata;  // mm_interconnect_0:credit_error_rx_0_s1_writedata -> credit_error_rx_0:writedata
	wire         mm_interconnect_0_data_en_to_w_s1_chipselect;      // mm_interconnect_0:data_en_to_w_s1_chipselect -> data_en_to_w:chipselect
	wire  [31:0] mm_interconnect_0_data_en_to_w_s1_readdata;        // data_en_to_w:readdata -> mm_interconnect_0:data_en_to_w_s1_readdata
	wire   [1:0] mm_interconnect_0_data_en_to_w_s1_address;         // mm_interconnect_0:data_en_to_w_s1_address -> data_en_to_w:address
	wire         mm_interconnect_0_data_en_to_w_s1_write;           // mm_interconnect_0:data_en_to_w_s1_write -> data_en_to_w:write_n
	wire  [31:0] mm_interconnect_0_data_en_to_w_s1_writedata;       // mm_interconnect_0:data_en_to_w_s1_writedata -> data_en_to_w:writedata
	wire         mm_interconnect_0_data_en_to_w_0_s1_chipselect;    // mm_interconnect_0:data_en_to_w_0_s1_chipselect -> data_en_to_w_0:chipselect
	wire  [31:0] mm_interconnect_0_data_en_to_w_0_s1_readdata;      // data_en_to_w_0:readdata -> mm_interconnect_0:data_en_to_w_0_s1_readdata
	wire   [1:0] mm_interconnect_0_data_en_to_w_0_s1_address;       // mm_interconnect_0:data_en_to_w_0_s1_address -> data_en_to_w_0:address
	wire         mm_interconnect_0_data_en_to_w_0_s1_write;         // mm_interconnect_0:data_en_to_w_0_s1_write -> data_en_to_w_0:write_n
	wire  [31:0] mm_interconnect_0_data_en_to_w_0_s1_writedata;     // mm_interconnect_0:data_en_to_w_0_s1_writedata -> data_en_to_w_0:writedata
	wire  [31:0] mm_interconnect_0_data_rx_r_s1_readdata;           // data_rx_r:readdata -> mm_interconnect_0:data_rx_r_s1_readdata
	wire   [1:0] mm_interconnect_0_data_rx_r_s1_address;            // mm_interconnect_0:data_rx_r_s1_address -> data_rx_r:address
	wire  [31:0] mm_interconnect_0_data_rx_r_0_s1_readdata;         // data_rx_r_0:readdata -> mm_interconnect_0:data_rx_r_0_s1_readdata
	wire   [1:0] mm_interconnect_0_data_rx_r_0_s1_address;          // mm_interconnect_0:data_rx_r_0_s1_address -> data_rx_r_0:address
	wire  [31:0] mm_interconnect_0_data_rx_ready_s1_readdata;       // data_rx_ready:readdata -> mm_interconnect_0:data_rx_ready_s1_readdata
	wire   [1:0] mm_interconnect_0_data_rx_ready_s1_address;        // mm_interconnect_0:data_rx_ready_s1_address -> data_rx_ready:address
	wire  [31:0] mm_interconnect_0_data_rx_ready_0_s1_readdata;     // data_rx_ready_0:readdata -> mm_interconnect_0:data_rx_ready_0_s1_readdata
	wire   [1:0] mm_interconnect_0_data_rx_ready_0_s1_address;      // mm_interconnect_0:data_rx_ready_0_s1_address -> data_rx_ready_0:address
	wire  [31:0] mm_interconnect_0_data_tx_ready_s1_readdata;       // data_tx_ready:readdata -> mm_interconnect_0:data_tx_ready_s1_readdata
	wire   [1:0] mm_interconnect_0_data_tx_ready_s1_address;        // mm_interconnect_0:data_tx_ready_s1_address -> data_tx_ready:address
	wire  [31:0] mm_interconnect_0_data_tx_ready_0_s1_readdata;     // data_tx_ready_0:readdata -> mm_interconnect_0:data_tx_ready_0_s1_readdata
	wire   [1:0] mm_interconnect_0_data_tx_ready_0_s1_address;      // mm_interconnect_0:data_tx_ready_0_s1_address -> data_tx_ready_0:address
	wire         mm_interconnect_0_data_tx_to_w_s1_chipselect;      // mm_interconnect_0:data_tx_to_w_s1_chipselect -> data_tx_to_w:chipselect
	wire  [31:0] mm_interconnect_0_data_tx_to_w_s1_readdata;        // data_tx_to_w:readdata -> mm_interconnect_0:data_tx_to_w_s1_readdata
	wire   [1:0] mm_interconnect_0_data_tx_to_w_s1_address;         // mm_interconnect_0:data_tx_to_w_s1_address -> data_tx_to_w:address
	wire         mm_interconnect_0_data_tx_to_w_s1_write;           // mm_interconnect_0:data_tx_to_w_s1_write -> data_tx_to_w:write_n
	wire  [31:0] mm_interconnect_0_data_tx_to_w_s1_writedata;       // mm_interconnect_0:data_tx_to_w_s1_writedata -> data_tx_to_w:writedata
	wire         mm_interconnect_0_data_tx_to_w_0_s1_chipselect;    // mm_interconnect_0:data_tx_to_w_0_s1_chipselect -> data_tx_to_w_0:chipselect
	wire  [31:0] mm_interconnect_0_data_tx_to_w_0_s1_readdata;      // data_tx_to_w_0:readdata -> mm_interconnect_0:data_tx_to_w_0_s1_readdata
	wire   [1:0] mm_interconnect_0_data_tx_to_w_0_s1_address;       // mm_interconnect_0:data_tx_to_w_0_s1_address -> data_tx_to_w_0:address
	wire         mm_interconnect_0_data_tx_to_w_0_s1_write;         // mm_interconnect_0:data_tx_to_w_0_s1_write -> data_tx_to_w_0:write_n
	wire  [31:0] mm_interconnect_0_data_tx_to_w_0_s1_writedata;     // mm_interconnect_0:data_tx_to_w_0_s1_writedata -> data_tx_to_w_0:writedata
	wire  [31:0] mm_interconnect_0_fsm_info_s1_readdata;            // fsm_info:readdata -> mm_interconnect_0:fsm_info_s1_readdata
	wire   [1:0] mm_interconnect_0_fsm_info_s1_address;             // mm_interconnect_0:fsm_info_s1_address -> fsm_info:address
	wire  [31:0] mm_interconnect_0_fsm_info_0_s1_readdata;          // fsm_info_0:readdata -> mm_interconnect_0:fsm_info_0_s1_readdata
	wire   [1:0] mm_interconnect_0_fsm_info_0_s1_address;           // mm_interconnect_0:fsm_info_0_s1_address -> fsm_info_0:address
	wire         mm_interconnect_0_link_disable_s1_chipselect;      // mm_interconnect_0:link_disable_s1_chipselect -> link_disable:chipselect
	wire  [31:0] mm_interconnect_0_link_disable_s1_readdata;        // link_disable:readdata -> mm_interconnect_0:link_disable_s1_readdata
	wire   [1:0] mm_interconnect_0_link_disable_s1_address;         // mm_interconnect_0:link_disable_s1_address -> link_disable:address
	wire         mm_interconnect_0_link_disable_s1_write;           // mm_interconnect_0:link_disable_s1_write -> link_disable:write_n
	wire  [31:0] mm_interconnect_0_link_disable_s1_writedata;       // mm_interconnect_0:link_disable_s1_writedata -> link_disable:writedata
	wire         mm_interconnect_0_link_disable_0_s1_chipselect;    // mm_interconnect_0:link_disable_0_s1_chipselect -> link_disable_0:chipselect
	wire  [31:0] mm_interconnect_0_link_disable_0_s1_readdata;      // link_disable_0:readdata -> mm_interconnect_0:link_disable_0_s1_readdata
	wire   [1:0] mm_interconnect_0_link_disable_0_s1_address;       // mm_interconnect_0:link_disable_0_s1_address -> link_disable_0:address
	wire         mm_interconnect_0_link_disable_0_s1_write;         // mm_interconnect_0:link_disable_0_s1_write -> link_disable_0:write_n
	wire  [31:0] mm_interconnect_0_link_disable_0_s1_writedata;     // mm_interconnect_0:link_disable_0_s1_writedata -> link_disable_0:writedata
	wire         mm_interconnect_0_link_start_s1_chipselect;        // mm_interconnect_0:link_start_s1_chipselect -> link_start:chipselect
	wire  [31:0] mm_interconnect_0_link_start_s1_readdata;          // link_start:readdata -> mm_interconnect_0:link_start_s1_readdata
	wire   [1:0] mm_interconnect_0_link_start_s1_address;           // mm_interconnect_0:link_start_s1_address -> link_start:address
	wire         mm_interconnect_0_link_start_s1_write;             // mm_interconnect_0:link_start_s1_write -> link_start:write_n
	wire  [31:0] mm_interconnect_0_link_start_s1_writedata;         // mm_interconnect_0:link_start_s1_writedata -> link_start:writedata
	wire         mm_interconnect_0_link_start_0_s1_chipselect;      // mm_interconnect_0:link_start_0_s1_chipselect -> link_start_0:chipselect
	wire  [31:0] mm_interconnect_0_link_start_0_s1_readdata;        // link_start_0:readdata -> mm_interconnect_0:link_start_0_s1_readdata
	wire   [1:0] mm_interconnect_0_link_start_0_s1_address;         // mm_interconnect_0:link_start_0_s1_address -> link_start_0:address
	wire         mm_interconnect_0_link_start_0_s1_write;           // mm_interconnect_0:link_start_0_s1_write -> link_start_0:write_n
	wire  [31:0] mm_interconnect_0_link_start_0_s1_writedata;       // mm_interconnect_0:link_start_0_s1_writedata -> link_start_0:writedata
	wire         mm_interconnect_0_send_fct_now_s1_chipselect;      // mm_interconnect_0:send_fct_now_s1_chipselect -> send_fct_now:chipselect
	wire  [31:0] mm_interconnect_0_send_fct_now_s1_readdata;        // send_fct_now:readdata -> mm_interconnect_0:send_fct_now_s1_readdata
	wire   [1:0] mm_interconnect_0_send_fct_now_s1_address;         // mm_interconnect_0:send_fct_now_s1_address -> send_fct_now:address
	wire         mm_interconnect_0_send_fct_now_s1_write;           // mm_interconnect_0:send_fct_now_s1_write -> send_fct_now:write_n
	wire  [31:0] mm_interconnect_0_send_fct_now_s1_writedata;       // mm_interconnect_0:send_fct_now_s1_writedata -> send_fct_now:writedata
	wire         mm_interconnect_0_send_fct_now_0_s1_chipselect;    // mm_interconnect_0:send_fct_now_0_s1_chipselect -> send_fct_now_0:chipselect
	wire  [31:0] mm_interconnect_0_send_fct_now_0_s1_readdata;      // send_fct_now_0:readdata -> mm_interconnect_0:send_fct_now_0_s1_readdata
	wire   [1:0] mm_interconnect_0_send_fct_now_0_s1_address;       // mm_interconnect_0:send_fct_now_0_s1_address -> send_fct_now_0:address
	wire         mm_interconnect_0_send_fct_now_0_s1_write;         // mm_interconnect_0:send_fct_now_0_s1_write -> send_fct_now_0:write_n
	wire  [31:0] mm_interconnect_0_send_fct_now_0_s1_writedata;     // mm_interconnect_0:send_fct_now_0_s1_writedata -> send_fct_now_0:writedata
	wire         mm_interconnect_0_timec_en_to_tx_s1_chipselect;    // mm_interconnect_0:timec_en_to_tx_s1_chipselect -> timec_en_to_tx:chipselect
	wire  [31:0] mm_interconnect_0_timec_en_to_tx_s1_readdata;      // timec_en_to_tx:readdata -> mm_interconnect_0:timec_en_to_tx_s1_readdata
	wire   [1:0] mm_interconnect_0_timec_en_to_tx_s1_address;       // mm_interconnect_0:timec_en_to_tx_s1_address -> timec_en_to_tx:address
	wire         mm_interconnect_0_timec_en_to_tx_s1_write;         // mm_interconnect_0:timec_en_to_tx_s1_write -> timec_en_to_tx:write_n
	wire  [31:0] mm_interconnect_0_timec_en_to_tx_s1_writedata;     // mm_interconnect_0:timec_en_to_tx_s1_writedata -> timec_en_to_tx:writedata
	wire         mm_interconnect_0_timec_en_to_tx_0_s1_chipselect;  // mm_interconnect_0:timec_en_to_tx_0_s1_chipselect -> timec_en_to_tx_0:chipselect
	wire  [31:0] mm_interconnect_0_timec_en_to_tx_0_s1_readdata;    // timec_en_to_tx_0:readdata -> mm_interconnect_0:timec_en_to_tx_0_s1_readdata
	wire   [1:0] mm_interconnect_0_timec_en_to_tx_0_s1_address;     // mm_interconnect_0:timec_en_to_tx_0_s1_address -> timec_en_to_tx_0:address
	wire         mm_interconnect_0_timec_en_to_tx_0_s1_write;       // mm_interconnect_0:timec_en_to_tx_0_s1_write -> timec_en_to_tx_0:write_n
	wire  [31:0] mm_interconnect_0_timec_en_to_tx_0_s1_writedata;   // mm_interconnect_0:timec_en_to_tx_0_s1_writedata -> timec_en_to_tx_0:writedata
	wire  [31:0] mm_interconnect_0_timec_rx_r_s1_readdata;          // timec_rx_r:readdata -> mm_interconnect_0:timec_rx_r_s1_readdata
	wire   [1:0] mm_interconnect_0_timec_rx_r_s1_address;           // mm_interconnect_0:timec_rx_r_s1_address -> timec_rx_r:address
	wire  [31:0] mm_interconnect_0_timec_rx_r_0_s1_readdata;        // timec_rx_r_0:readdata -> mm_interconnect_0:timec_rx_r_0_s1_readdata
	wire   [1:0] mm_interconnect_0_timec_rx_r_0_s1_address;         // mm_interconnect_0:timec_rx_r_0_s1_address -> timec_rx_r_0:address
	wire  [31:0] mm_interconnect_0_timec_rx_ready_s1_readdata;      // timec_rx_ready:readdata -> mm_interconnect_0:timec_rx_ready_s1_readdata
	wire   [1:0] mm_interconnect_0_timec_rx_ready_s1_address;       // mm_interconnect_0:timec_rx_ready_s1_address -> timec_rx_ready:address
	wire  [31:0] mm_interconnect_0_timec_rx_ready_0_s1_readdata;    // timec_rx_ready_0:readdata -> mm_interconnect_0:timec_rx_ready_0_s1_readdata
	wire   [1:0] mm_interconnect_0_timec_rx_ready_0_s1_address;     // mm_interconnect_0:timec_rx_ready_0_s1_address -> timec_rx_ready_0:address
	wire  [31:0] mm_interconnect_0_timec_tx_ready_s1_readdata;      // timec_tx_ready:readdata -> mm_interconnect_0:timec_tx_ready_s1_readdata
	wire   [1:0] mm_interconnect_0_timec_tx_ready_s1_address;       // mm_interconnect_0:timec_tx_ready_s1_address -> timec_tx_ready:address
	wire  [31:0] mm_interconnect_0_timec_tx_ready_0_s1_readdata;    // timec_tx_ready_0:readdata -> mm_interconnect_0:timec_tx_ready_0_s1_readdata
	wire   [1:0] mm_interconnect_0_timec_tx_ready_0_s1_address;     // mm_interconnect_0:timec_tx_ready_0_s1_address -> timec_tx_ready_0:address
	wire         mm_interconnect_0_timec_tx_to_w_s1_chipselect;     // mm_interconnect_0:timec_tx_to_w_s1_chipselect -> timec_tx_to_w:chipselect
	wire  [31:0] mm_interconnect_0_timec_tx_to_w_s1_readdata;       // timec_tx_to_w:readdata -> mm_interconnect_0:timec_tx_to_w_s1_readdata
	wire   [1:0] mm_interconnect_0_timec_tx_to_w_s1_address;        // mm_interconnect_0:timec_tx_to_w_s1_address -> timec_tx_to_w:address
	wire         mm_interconnect_0_timec_tx_to_w_s1_write;          // mm_interconnect_0:timec_tx_to_w_s1_write -> timec_tx_to_w:write_n
	wire  [31:0] mm_interconnect_0_timec_tx_to_w_s1_writedata;      // mm_interconnect_0:timec_tx_to_w_s1_writedata -> timec_tx_to_w:writedata
	wire         mm_interconnect_0_timec_tx_to_w_0_s1_chipselect;   // mm_interconnect_0:timec_tx_to_w_0_s1_chipselect -> timec_tx_to_w_0:chipselect
	wire  [31:0] mm_interconnect_0_timec_tx_to_w_0_s1_readdata;     // timec_tx_to_w_0:readdata -> mm_interconnect_0:timec_tx_to_w_0_s1_readdata
	wire   [1:0] mm_interconnect_0_timec_tx_to_w_0_s1_address;      // mm_interconnect_0:timec_tx_to_w_0_s1_address -> timec_tx_to_w_0:address
	wire         mm_interconnect_0_timec_tx_to_w_0_s1_write;        // mm_interconnect_0:timec_tx_to_w_0_s1_write -> timec_tx_to_w_0:write_n
	wire  [31:0] mm_interconnect_0_timec_tx_to_w_0_s1_writedata;    // mm_interconnect_0:timec_tx_to_w_0_s1_writedata -> timec_tx_to_w_0:writedata
	wire         rst_controller_reset_out_reset;                    // rst_controller:reset_out -> [MONITOR_A:reset_n, MONITOR_B:reset_n, auto_start:reset_n, auto_start_0:reset_n, clock_sel:reset_n, credit_error_rx:reset_n, credit_error_rx_0:reset_n, data_en_to_w:reset_n, data_en_to_w_0:reset_n, data_rx_r:reset_n, data_rx_r_0:reset_n, data_rx_ready:reset_n, data_rx_ready_0:reset_n, data_tx_ready:reset_n, data_tx_ready_0:reset_n, data_tx_to_w:reset_n, data_tx_to_w_0:reset_n, fsm_info:reset_n, fsm_info_0:reset_n, led_fpga:reset_n, link_disable:reset_n, link_disable_0:reset_n, link_start:reset_n, link_start_0:reset_n, mm_interconnect_0:led_fpga_reset_reset_bridge_in_reset_reset, send_fct_now:reset_n, send_fct_now_0:reset_n, timec_en_to_tx:reset_n, timec_en_to_tx_0:reset_n, timec_rx_r:reset_n, timec_rx_r_0:reset_n, timec_rx_ready:reset_n, timec_rx_ready_0:reset_n, timec_tx_ready:reset_n, timec_tx_ready_0:reset_n, timec_tx_to_w:reset_n, timec_tx_to_w_0:reset_n]
	wire         rst_controller_001_reset_out_reset;                // rst_controller_001:reset_out -> mm_interconnect_0:hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset
	wire         hps_0_h2f_reset_reset;                             // hps_0:h2f_rst_n -> rst_controller_001:reset_in0

	spw_ulight_nofifo_MONITOR_A monitor_a (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address  (mm_interconnect_0_monitor_a_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_monitor_a_s1_readdata), //                    .readdata
		.in_port  (monitor_a_external_connection_export)     // external_connection.export
	);

	spw_ulight_nofifo_MONITOR_A monitor_b (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address  (mm_interconnect_0_monitor_b_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_monitor_b_s1_readdata), //                    .readdata
		.in_port  (monitor_b_external_connection_export)     // external_connection.export
	);

	spw_ulight_nofifo_auto_start auto_start (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_auto_start_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_auto_start_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_auto_start_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_auto_start_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_auto_start_s1_readdata),   //                    .readdata
		.out_port   (auto_start_external_connection_export)       // external_connection.export
	);

	spw_ulight_nofifo_auto_start auto_start_0 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_auto_start_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_auto_start_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_auto_start_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_auto_start_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_auto_start_0_s1_readdata),   //                    .readdata
		.out_port   (auto_start_0_external_connection_export)       // external_connection.export
	);

	spw_ulight_nofifo_clock_sel clock_sel (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_clock_sel_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_clock_sel_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_clock_sel_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_clock_sel_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_clock_sel_s1_readdata),   //                    .readdata
		.out_port   (clock_sel_external_connection_export)       // external_connection.export
	);

	spw_ulight_nofifo_auto_start credit_error_rx (
		.clk        (clk_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_credit_error_rx_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_credit_error_rx_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_credit_error_rx_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_credit_error_rx_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_credit_error_rx_s1_readdata),   //                    .readdata
		.out_port   (credit_error_rx_external_connection_export)       // external_connection.export
	);

	spw_ulight_nofifo_auto_start credit_error_rx_0 (
		.clk        (clk_clk),                                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (mm_interconnect_0_credit_error_rx_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_credit_error_rx_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_credit_error_rx_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_credit_error_rx_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_credit_error_rx_0_s1_readdata),   //                    .readdata
		.out_port   (credit_error_rx_0_external_connection_export)       // external_connection.export
	);

	spw_ulight_nofifo_auto_start data_en_to_w (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_data_en_to_w_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_data_en_to_w_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_data_en_to_w_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_data_en_to_w_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_data_en_to_w_s1_readdata),   //                    .readdata
		.out_port   (data_en_to_w_external_connection_export)       // external_connection.export
	);

	spw_ulight_nofifo_auto_start data_en_to_w_0 (
		.clk        (clk_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_data_en_to_w_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_data_en_to_w_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_data_en_to_w_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_data_en_to_w_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_data_en_to_w_0_s1_readdata),   //                    .readdata
		.out_port   (data_en_to_w_0_external_connection_export)       // external_connection.export
	);

	spw_ulight_nofifo_data_rx_r data_rx_r (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address  (mm_interconnect_0_data_rx_r_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_data_rx_r_s1_readdata), //                    .readdata
		.in_port  (data_rx_r_external_connection_export)     // external_connection.export
	);

	spw_ulight_nofifo_data_rx_r data_rx_r_0 (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_0_data_rx_r_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_data_rx_r_0_s1_readdata), //                    .readdata
		.in_port  (data_rx_r_0_external_connection_export)     // external_connection.export
	);

	spw_ulight_nofifo_data_rx_ready data_rx_ready (
		.clk      (clk_clk),                                     //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address  (mm_interconnect_0_data_rx_ready_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_data_rx_ready_s1_readdata), //                    .readdata
		.in_port  (data_rx_ready_external_connection_export)     // external_connection.export
	);

	spw_ulight_nofifo_data_rx_ready data_rx_ready_0 (
		.clk      (clk_clk),                                       //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address  (mm_interconnect_0_data_rx_ready_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_data_rx_ready_0_s1_readdata), //                    .readdata
		.in_port  (data_rx_ready_0_external_connection_export)     // external_connection.export
	);

	spw_ulight_nofifo_data_rx_ready data_tx_ready (
		.clk      (clk_clk),                                     //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address  (mm_interconnect_0_data_tx_ready_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_data_tx_ready_s1_readdata), //                    .readdata
		.in_port  (data_tx_ready_external_connection_export)     // external_connection.export
	);

	spw_ulight_nofifo_data_rx_ready data_tx_ready_0 (
		.clk      (clk_clk),                                       //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address  (mm_interconnect_0_data_tx_ready_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_data_tx_ready_0_s1_readdata), //                    .readdata
		.in_port  (data_tx_ready_0_external_connection_export)     // external_connection.export
	);

	spw_ulight_nofifo_data_tx_to_w data_tx_to_w (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_data_tx_to_w_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_data_tx_to_w_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_data_tx_to_w_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_data_tx_to_w_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_data_tx_to_w_s1_readdata),   //                    .readdata
		.out_port   (data_tx_to_w_external_connection_export)       // external_connection.export
	);

	spw_ulight_nofifo_data_tx_to_w data_tx_to_w_0 (
		.clk        (clk_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_data_tx_to_w_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_data_tx_to_w_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_data_tx_to_w_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_data_tx_to_w_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_data_tx_to_w_0_s1_readdata),   //                    .readdata
		.out_port   (data_tx_to_w_0_external_connection_export)       // external_connection.export
	);

	spw_ulight_nofifo_fsm_info fsm_info (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_fsm_info_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_fsm_info_s1_readdata), //                    .readdata
		.in_port  (fsm_info_external_connection_export)     // external_connection.export
	);

	spw_ulight_nofifo_fsm_info fsm_info_0 (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_fsm_info_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_fsm_info_0_s1_readdata), //                    .readdata
		.in_port  (fsm_info_0_external_connection_export)     // external_connection.export
	);

	spw_ulight_nofifo_hps_0 #(
		.F2S_Width (0),
		.S2F_Width (1)
	) hps_0 (
		.mem_a          (),                             //            memory.mem_a
		.mem_ba         (),                             //                  .mem_ba
		.mem_ck         (),                             //                  .mem_ck
		.mem_ck_n       (),                             //                  .mem_ck_n
		.mem_cke        (),                             //                  .mem_cke
		.mem_cs_n       (),                             //                  .mem_cs_n
		.mem_ras_n      (),                             //                  .mem_ras_n
		.mem_cas_n      (),                             //                  .mem_cas_n
		.mem_we_n       (),                             //                  .mem_we_n
		.mem_reset_n    (),                             //                  .mem_reset_n
		.mem_dq         (),                             //                  .mem_dq
		.mem_dqs        (),                             //                  .mem_dqs
		.mem_dqs_n      (),                             //                  .mem_dqs_n
		.mem_odt        (),                             //                  .mem_odt
		.mem_dm         (),                             //                  .mem_dm
		.oct_rzqin      (),                             //                  .oct_rzqin
		.h2f_rst_n      (hps_0_h2f_reset_reset),        //         h2f_reset.reset_n
		.h2f_axi_clk    (clk_clk),                      //     h2f_axi_clock.clk
		.h2f_AWID       (hps_0_h2f_axi_master_awid),    //    h2f_axi_master.awid
		.h2f_AWADDR     (hps_0_h2f_axi_master_awaddr),  //                  .awaddr
		.h2f_AWLEN      (hps_0_h2f_axi_master_awlen),   //                  .awlen
		.h2f_AWSIZE     (hps_0_h2f_axi_master_awsize),  //                  .awsize
		.h2f_AWBURST    (hps_0_h2f_axi_master_awburst), //                  .awburst
		.h2f_AWLOCK     (hps_0_h2f_axi_master_awlock),  //                  .awlock
		.h2f_AWCACHE    (hps_0_h2f_axi_master_awcache), //                  .awcache
		.h2f_AWPROT     (hps_0_h2f_axi_master_awprot),  //                  .awprot
		.h2f_AWVALID    (hps_0_h2f_axi_master_awvalid), //                  .awvalid
		.h2f_AWREADY    (hps_0_h2f_axi_master_awready), //                  .awready
		.h2f_WID        (hps_0_h2f_axi_master_wid),     //                  .wid
		.h2f_WDATA      (hps_0_h2f_axi_master_wdata),   //                  .wdata
		.h2f_WSTRB      (hps_0_h2f_axi_master_wstrb),   //                  .wstrb
		.h2f_WLAST      (hps_0_h2f_axi_master_wlast),   //                  .wlast
		.h2f_WVALID     (hps_0_h2f_axi_master_wvalid),  //                  .wvalid
		.h2f_WREADY     (hps_0_h2f_axi_master_wready),  //                  .wready
		.h2f_BID        (hps_0_h2f_axi_master_bid),     //                  .bid
		.h2f_BRESP      (hps_0_h2f_axi_master_bresp),   //                  .bresp
		.h2f_BVALID     (hps_0_h2f_axi_master_bvalid),  //                  .bvalid
		.h2f_BREADY     (hps_0_h2f_axi_master_bready),  //                  .bready
		.h2f_ARID       (hps_0_h2f_axi_master_arid),    //                  .arid
		.h2f_ARADDR     (hps_0_h2f_axi_master_araddr),  //                  .araddr
		.h2f_ARLEN      (hps_0_h2f_axi_master_arlen),   //                  .arlen
		.h2f_ARSIZE     (hps_0_h2f_axi_master_arsize),  //                  .arsize
		.h2f_ARBURST    (hps_0_h2f_axi_master_arburst), //                  .arburst
		.h2f_ARLOCK     (hps_0_h2f_axi_master_arlock),  //                  .arlock
		.h2f_ARCACHE    (hps_0_h2f_axi_master_arcache), //                  .arcache
		.h2f_ARPROT     (hps_0_h2f_axi_master_arprot),  //                  .arprot
		.h2f_ARVALID    (hps_0_h2f_axi_master_arvalid), //                  .arvalid
		.h2f_ARREADY    (hps_0_h2f_axi_master_arready), //                  .arready
		.h2f_RID        (hps_0_h2f_axi_master_rid),     //                  .rid
		.h2f_RDATA      (hps_0_h2f_axi_master_rdata),   //                  .rdata
		.h2f_RRESP      (hps_0_h2f_axi_master_rresp),   //                  .rresp
		.h2f_RLAST      (hps_0_h2f_axi_master_rlast),   //                  .rlast
		.h2f_RVALID     (hps_0_h2f_axi_master_rvalid),  //                  .rvalid
		.h2f_RREADY     (hps_0_h2f_axi_master_rready),  //                  .rready
		.h2f_lw_axi_clk (clk_clk),                      //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID    (),                             // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR  (),                             //                  .awaddr
		.h2f_lw_AWLEN   (),                             //                  .awlen
		.h2f_lw_AWSIZE  (),                             //                  .awsize
		.h2f_lw_AWBURST (),                             //                  .awburst
		.h2f_lw_AWLOCK  (),                             //                  .awlock
		.h2f_lw_AWCACHE (),                             //                  .awcache
		.h2f_lw_AWPROT  (),                             //                  .awprot
		.h2f_lw_AWVALID (),                             //                  .awvalid
		.h2f_lw_AWREADY (),                             //                  .awready
		.h2f_lw_WID     (),                             //                  .wid
		.h2f_lw_WDATA   (),                             //                  .wdata
		.h2f_lw_WSTRB   (),                             //                  .wstrb
		.h2f_lw_WLAST   (),                             //                  .wlast
		.h2f_lw_WVALID  (),                             //                  .wvalid
		.h2f_lw_WREADY  (),                             //                  .wready
		.h2f_lw_BID     (),                             //                  .bid
		.h2f_lw_BRESP   (),                             //                  .bresp
		.h2f_lw_BVALID  (),                             //                  .bvalid
		.h2f_lw_BREADY  (),                             //                  .bready
		.h2f_lw_ARID    (),                             //                  .arid
		.h2f_lw_ARADDR  (),                             //                  .araddr
		.h2f_lw_ARLEN   (),                             //                  .arlen
		.h2f_lw_ARSIZE  (),                             //                  .arsize
		.h2f_lw_ARBURST (),                             //                  .arburst
		.h2f_lw_ARLOCK  (),                             //                  .arlock
		.h2f_lw_ARCACHE (),                             //                  .arcache
		.h2f_lw_ARPROT  (),                             //                  .arprot
		.h2f_lw_ARVALID (),                             //                  .arvalid
		.h2f_lw_ARREADY (),                             //                  .arready
		.h2f_lw_RID     (),                             //                  .rid
		.h2f_lw_RDATA   (),                             //                  .rdata
		.h2f_lw_RRESP   (),                             //                  .rresp
		.h2f_lw_RLAST   (),                             //                  .rlast
		.h2f_lw_RVALID  (),                             //                  .rvalid
		.h2f_lw_RREADY  ()                              //                  .rready
	);

	spw_ulight_nofifo_led_fpga led_fpga (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_led_fpga_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_fpga_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_fpga_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_fpga_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_fpga_s1_readdata),   //                    .readdata
		.out_port   (led_fpga_external_connection_export)       // external_connection.export
	);

	spw_ulight_nofifo_auto_start link_disable (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_link_disable_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_link_disable_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_link_disable_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_link_disable_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_link_disable_s1_readdata),   //                    .readdata
		.out_port   (link_disable_external_connection_export)       // external_connection.export
	);

	spw_ulight_nofifo_auto_start link_disable_0 (
		.clk        (clk_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_link_disable_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_link_disable_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_link_disable_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_link_disable_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_link_disable_0_s1_readdata),   //                    .readdata
		.out_port   (link_disable_0_external_connection_export)       // external_connection.export
	);

	spw_ulight_nofifo_auto_start link_start (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_link_start_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_link_start_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_link_start_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_link_start_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_link_start_s1_readdata),   //                    .readdata
		.out_port   (link_start_external_connection_export)       // external_connection.export
	);

	spw_ulight_nofifo_auto_start link_start_0 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_link_start_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_link_start_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_link_start_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_link_start_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_link_start_0_s1_readdata),   //                    .readdata
		.out_port   (link_start_0_external_connection_export)       // external_connection.export
	);

	spw_ulight_nofifo_pll_tx pll_tx (
		.refclk   (clk_clk),              //  refclk.clk
		.rst      (~reset_reset_n),       //   reset.reset
		.outclk_0 (pll_tx_outclk0_clk),   // outclk0.clk
		.outclk_1 (pll_tx_outclk1_clk),   // outclk1.clk
		.outclk_2 (pll_tx_outclk2_clk),   // outclk2.clk
		.outclk_3 (pll_tx_outclk3_clk),   // outclk3.clk
		.outclk_4 (pll_tx_outclk4_clk),   // outclk4.clk
		.locked   (pll_tx_locked_export), //  locked.export
		.refclk1  ()                      // refclk1.refclk1
	);

	spw_ulight_nofifo_auto_start send_fct_now (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_send_fct_now_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_send_fct_now_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_send_fct_now_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_send_fct_now_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_send_fct_now_s1_readdata),   //                    .readdata
		.out_port   (send_fct_now_external_connection_export)       // external_connection.export
	);

	spw_ulight_nofifo_auto_start send_fct_now_0 (
		.clk        (clk_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_send_fct_now_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_send_fct_now_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_send_fct_now_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_send_fct_now_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_send_fct_now_0_s1_readdata),   //                    .readdata
		.out_port   (send_fct_now_0_external_connection_export)       // external_connection.export
	);

	spw_ulight_nofifo_auto_start timec_en_to_tx (
		.clk        (clk_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_timec_en_to_tx_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_timec_en_to_tx_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_timec_en_to_tx_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_timec_en_to_tx_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_timec_en_to_tx_s1_readdata),   //                    .readdata
		.out_port   (timec_en_to_tx_external_connection_export)       // external_connection.export
	);

	spw_ulight_nofifo_auto_start timec_en_to_tx_0 (
		.clk        (clk_clk),                                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (mm_interconnect_0_timec_en_to_tx_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_timec_en_to_tx_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_timec_en_to_tx_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_timec_en_to_tx_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_timec_en_to_tx_0_s1_readdata),   //                    .readdata
		.out_port   (timec_en_to_tx_0_external_connection_export)       // external_connection.export
	);

	spw_ulight_nofifo_timec_rx_r timec_rx_r (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_timec_rx_r_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_timec_rx_r_s1_readdata), //                    .readdata
		.in_port  (timec_rx_r_external_connection_export)     // external_connection.export
	);

	spw_ulight_nofifo_timec_rx_r timec_rx_r_0 (
		.clk      (clk_clk),                                    //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_0_timec_rx_r_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_timec_rx_r_0_s1_readdata), //                    .readdata
		.in_port  (timec_rx_r_0_external_connection_export)     // external_connection.export
	);

	spw_ulight_nofifo_data_rx_ready timec_rx_ready (
		.clk      (clk_clk),                                      //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address  (mm_interconnect_0_timec_rx_ready_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_timec_rx_ready_s1_readdata), //                    .readdata
		.in_port  (timec_rx_ready_external_connection_export)     // external_connection.export
	);

	spw_ulight_nofifo_data_rx_ready timec_rx_ready_0 (
		.clk      (clk_clk),                                        //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address  (mm_interconnect_0_timec_rx_ready_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_timec_rx_ready_0_s1_readdata), //                    .readdata
		.in_port  (timec_rx_ready_0_external_connection_export)     // external_connection.export
	);

	spw_ulight_nofifo_data_rx_ready timec_tx_ready (
		.clk      (clk_clk),                                      //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address  (mm_interconnect_0_timec_tx_ready_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_timec_tx_ready_s1_readdata), //                    .readdata
		.in_port  (timec_tx_ready_external_connection_export)     // external_connection.export
	);

	spw_ulight_nofifo_data_rx_ready timec_tx_ready_0 (
		.clk      (clk_clk),                                        //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address  (mm_interconnect_0_timec_tx_ready_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_timec_tx_ready_0_s1_readdata), //                    .readdata
		.in_port  (timec_tx_ready_0_external_connection_export)     // external_connection.export
	);

	spw_ulight_nofifo_timec_tx_to_w timec_tx_to_w (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_timec_tx_to_w_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_timec_tx_to_w_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_timec_tx_to_w_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_timec_tx_to_w_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_timec_tx_to_w_s1_readdata),   //                    .readdata
		.out_port   (timec_tx_to_w_external_connection_export)       // external_connection.export
	);

	spw_ulight_nofifo_timec_tx_to_w timec_tx_to_w_0 (
		.clk        (clk_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_timec_tx_to_w_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_timec_tx_to_w_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_timec_tx_to_w_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_timec_tx_to_w_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_timec_tx_to_w_0_s1_readdata),   //                    .readdata
		.out_port   (timec_tx_to_w_0_external_connection_export)       // external_connection.export
	);

	spw_ulight_nofifo_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_h2f_axi_master_awid                                        (hps_0_h2f_axi_master_awid),                         //                                       hps_0_h2f_axi_master.awid
		.hps_0_h2f_axi_master_awaddr                                      (hps_0_h2f_axi_master_awaddr),                       //                                                           .awaddr
		.hps_0_h2f_axi_master_awlen                                       (hps_0_h2f_axi_master_awlen),                        //                                                           .awlen
		.hps_0_h2f_axi_master_awsize                                      (hps_0_h2f_axi_master_awsize),                       //                                                           .awsize
		.hps_0_h2f_axi_master_awburst                                     (hps_0_h2f_axi_master_awburst),                      //                                                           .awburst
		.hps_0_h2f_axi_master_awlock                                      (hps_0_h2f_axi_master_awlock),                       //                                                           .awlock
		.hps_0_h2f_axi_master_awcache                                     (hps_0_h2f_axi_master_awcache),                      //                                                           .awcache
		.hps_0_h2f_axi_master_awprot                                      (hps_0_h2f_axi_master_awprot),                       //                                                           .awprot
		.hps_0_h2f_axi_master_awvalid                                     (hps_0_h2f_axi_master_awvalid),                      //                                                           .awvalid
		.hps_0_h2f_axi_master_awready                                     (hps_0_h2f_axi_master_awready),                      //                                                           .awready
		.hps_0_h2f_axi_master_wid                                         (hps_0_h2f_axi_master_wid),                          //                                                           .wid
		.hps_0_h2f_axi_master_wdata                                       (hps_0_h2f_axi_master_wdata),                        //                                                           .wdata
		.hps_0_h2f_axi_master_wstrb                                       (hps_0_h2f_axi_master_wstrb),                        //                                                           .wstrb
		.hps_0_h2f_axi_master_wlast                                       (hps_0_h2f_axi_master_wlast),                        //                                                           .wlast
		.hps_0_h2f_axi_master_wvalid                                      (hps_0_h2f_axi_master_wvalid),                       //                                                           .wvalid
		.hps_0_h2f_axi_master_wready                                      (hps_0_h2f_axi_master_wready),                       //                                                           .wready
		.hps_0_h2f_axi_master_bid                                         (hps_0_h2f_axi_master_bid),                          //                                                           .bid
		.hps_0_h2f_axi_master_bresp                                       (hps_0_h2f_axi_master_bresp),                        //                                                           .bresp
		.hps_0_h2f_axi_master_bvalid                                      (hps_0_h2f_axi_master_bvalid),                       //                                                           .bvalid
		.hps_0_h2f_axi_master_bready                                      (hps_0_h2f_axi_master_bready),                       //                                                           .bready
		.hps_0_h2f_axi_master_arid                                        (hps_0_h2f_axi_master_arid),                         //                                                           .arid
		.hps_0_h2f_axi_master_araddr                                      (hps_0_h2f_axi_master_araddr),                       //                                                           .araddr
		.hps_0_h2f_axi_master_arlen                                       (hps_0_h2f_axi_master_arlen),                        //                                                           .arlen
		.hps_0_h2f_axi_master_arsize                                      (hps_0_h2f_axi_master_arsize),                       //                                                           .arsize
		.hps_0_h2f_axi_master_arburst                                     (hps_0_h2f_axi_master_arburst),                      //                                                           .arburst
		.hps_0_h2f_axi_master_arlock                                      (hps_0_h2f_axi_master_arlock),                       //                                                           .arlock
		.hps_0_h2f_axi_master_arcache                                     (hps_0_h2f_axi_master_arcache),                      //                                                           .arcache
		.hps_0_h2f_axi_master_arprot                                      (hps_0_h2f_axi_master_arprot),                       //                                                           .arprot
		.hps_0_h2f_axi_master_arvalid                                     (hps_0_h2f_axi_master_arvalid),                      //                                                           .arvalid
		.hps_0_h2f_axi_master_arready                                     (hps_0_h2f_axi_master_arready),                      //                                                           .arready
		.hps_0_h2f_axi_master_rid                                         (hps_0_h2f_axi_master_rid),                          //                                                           .rid
		.hps_0_h2f_axi_master_rdata                                       (hps_0_h2f_axi_master_rdata),                        //                                                           .rdata
		.hps_0_h2f_axi_master_rresp                                       (hps_0_h2f_axi_master_rresp),                        //                                                           .rresp
		.hps_0_h2f_axi_master_rlast                                       (hps_0_h2f_axi_master_rlast),                        //                                                           .rlast
		.hps_0_h2f_axi_master_rvalid                                      (hps_0_h2f_axi_master_rvalid),                       //                                                           .rvalid
		.hps_0_h2f_axi_master_rready                                      (hps_0_h2f_axi_master_rready),                       //                                                           .rready
		.clk_0_clk_clk                                                    (clk_clk),                                           //                                                  clk_0_clk.clk
		.hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                // hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.led_fpga_reset_reset_bridge_in_reset_reset                       (rst_controller_reset_out_reset),                    //                       led_fpga_reset_reset_bridge_in_reset.reset
		.auto_start_s1_address                                            (mm_interconnect_0_auto_start_s1_address),           //                                              auto_start_s1.address
		.auto_start_s1_write                                              (mm_interconnect_0_auto_start_s1_write),             //                                                           .write
		.auto_start_s1_readdata                                           (mm_interconnect_0_auto_start_s1_readdata),          //                                                           .readdata
		.auto_start_s1_writedata                                          (mm_interconnect_0_auto_start_s1_writedata),         //                                                           .writedata
		.auto_start_s1_chipselect                                         (mm_interconnect_0_auto_start_s1_chipselect),        //                                                           .chipselect
		.auto_start_0_s1_address                                          (mm_interconnect_0_auto_start_0_s1_address),         //                                            auto_start_0_s1.address
		.auto_start_0_s1_write                                            (mm_interconnect_0_auto_start_0_s1_write),           //                                                           .write
		.auto_start_0_s1_readdata                                         (mm_interconnect_0_auto_start_0_s1_readdata),        //                                                           .readdata
		.auto_start_0_s1_writedata                                        (mm_interconnect_0_auto_start_0_s1_writedata),       //                                                           .writedata
		.auto_start_0_s1_chipselect                                       (mm_interconnect_0_auto_start_0_s1_chipselect),      //                                                           .chipselect
		.clock_sel_s1_address                                             (mm_interconnect_0_clock_sel_s1_address),            //                                               clock_sel_s1.address
		.clock_sel_s1_write                                               (mm_interconnect_0_clock_sel_s1_write),              //                                                           .write
		.clock_sel_s1_readdata                                            (mm_interconnect_0_clock_sel_s1_readdata),           //                                                           .readdata
		.clock_sel_s1_writedata                                           (mm_interconnect_0_clock_sel_s1_writedata),          //                                                           .writedata
		.clock_sel_s1_chipselect                                          (mm_interconnect_0_clock_sel_s1_chipselect),         //                                                           .chipselect
		.credit_error_rx_s1_address                                       (mm_interconnect_0_credit_error_rx_s1_address),      //                                         credit_error_rx_s1.address
		.credit_error_rx_s1_write                                         (mm_interconnect_0_credit_error_rx_s1_write),        //                                                           .write
		.credit_error_rx_s1_readdata                                      (mm_interconnect_0_credit_error_rx_s1_readdata),     //                                                           .readdata
		.credit_error_rx_s1_writedata                                     (mm_interconnect_0_credit_error_rx_s1_writedata),    //                                                           .writedata
		.credit_error_rx_s1_chipselect                                    (mm_interconnect_0_credit_error_rx_s1_chipselect),   //                                                           .chipselect
		.credit_error_rx_0_s1_address                                     (mm_interconnect_0_credit_error_rx_0_s1_address),    //                                       credit_error_rx_0_s1.address
		.credit_error_rx_0_s1_write                                       (mm_interconnect_0_credit_error_rx_0_s1_write),      //                                                           .write
		.credit_error_rx_0_s1_readdata                                    (mm_interconnect_0_credit_error_rx_0_s1_readdata),   //                                                           .readdata
		.credit_error_rx_0_s1_writedata                                   (mm_interconnect_0_credit_error_rx_0_s1_writedata),  //                                                           .writedata
		.credit_error_rx_0_s1_chipselect                                  (mm_interconnect_0_credit_error_rx_0_s1_chipselect), //                                                           .chipselect
		.data_en_to_w_s1_address                                          (mm_interconnect_0_data_en_to_w_s1_address),         //                                            data_en_to_w_s1.address
		.data_en_to_w_s1_write                                            (mm_interconnect_0_data_en_to_w_s1_write),           //                                                           .write
		.data_en_to_w_s1_readdata                                         (mm_interconnect_0_data_en_to_w_s1_readdata),        //                                                           .readdata
		.data_en_to_w_s1_writedata                                        (mm_interconnect_0_data_en_to_w_s1_writedata),       //                                                           .writedata
		.data_en_to_w_s1_chipselect                                       (mm_interconnect_0_data_en_to_w_s1_chipselect),      //                                                           .chipselect
		.data_en_to_w_0_s1_address                                        (mm_interconnect_0_data_en_to_w_0_s1_address),       //                                          data_en_to_w_0_s1.address
		.data_en_to_w_0_s1_write                                          (mm_interconnect_0_data_en_to_w_0_s1_write),         //                                                           .write
		.data_en_to_w_0_s1_readdata                                       (mm_interconnect_0_data_en_to_w_0_s1_readdata),      //                                                           .readdata
		.data_en_to_w_0_s1_writedata                                      (mm_interconnect_0_data_en_to_w_0_s1_writedata),     //                                                           .writedata
		.data_en_to_w_0_s1_chipselect                                     (mm_interconnect_0_data_en_to_w_0_s1_chipselect),    //                                                           .chipselect
		.data_rx_r_s1_address                                             (mm_interconnect_0_data_rx_r_s1_address),            //                                               data_rx_r_s1.address
		.data_rx_r_s1_readdata                                            (mm_interconnect_0_data_rx_r_s1_readdata),           //                                                           .readdata
		.data_rx_r_0_s1_address                                           (mm_interconnect_0_data_rx_r_0_s1_address),          //                                             data_rx_r_0_s1.address
		.data_rx_r_0_s1_readdata                                          (mm_interconnect_0_data_rx_r_0_s1_readdata),         //                                                           .readdata
		.data_rx_ready_s1_address                                         (mm_interconnect_0_data_rx_ready_s1_address),        //                                           data_rx_ready_s1.address
		.data_rx_ready_s1_readdata                                        (mm_interconnect_0_data_rx_ready_s1_readdata),       //                                                           .readdata
		.data_rx_ready_0_s1_address                                       (mm_interconnect_0_data_rx_ready_0_s1_address),      //                                         data_rx_ready_0_s1.address
		.data_rx_ready_0_s1_readdata                                      (mm_interconnect_0_data_rx_ready_0_s1_readdata),     //                                                           .readdata
		.data_tx_ready_s1_address                                         (mm_interconnect_0_data_tx_ready_s1_address),        //                                           data_tx_ready_s1.address
		.data_tx_ready_s1_readdata                                        (mm_interconnect_0_data_tx_ready_s1_readdata),       //                                                           .readdata
		.data_tx_ready_0_s1_address                                       (mm_interconnect_0_data_tx_ready_0_s1_address),      //                                         data_tx_ready_0_s1.address
		.data_tx_ready_0_s1_readdata                                      (mm_interconnect_0_data_tx_ready_0_s1_readdata),     //                                                           .readdata
		.data_tx_to_w_s1_address                                          (mm_interconnect_0_data_tx_to_w_s1_address),         //                                            data_tx_to_w_s1.address
		.data_tx_to_w_s1_write                                            (mm_interconnect_0_data_tx_to_w_s1_write),           //                                                           .write
		.data_tx_to_w_s1_readdata                                         (mm_interconnect_0_data_tx_to_w_s1_readdata),        //                                                           .readdata
		.data_tx_to_w_s1_writedata                                        (mm_interconnect_0_data_tx_to_w_s1_writedata),       //                                                           .writedata
		.data_tx_to_w_s1_chipselect                                       (mm_interconnect_0_data_tx_to_w_s1_chipselect),      //                                                           .chipselect
		.data_tx_to_w_0_s1_address                                        (mm_interconnect_0_data_tx_to_w_0_s1_address),       //                                          data_tx_to_w_0_s1.address
		.data_tx_to_w_0_s1_write                                          (mm_interconnect_0_data_tx_to_w_0_s1_write),         //                                                           .write
		.data_tx_to_w_0_s1_readdata                                       (mm_interconnect_0_data_tx_to_w_0_s1_readdata),      //                                                           .readdata
		.data_tx_to_w_0_s1_writedata                                      (mm_interconnect_0_data_tx_to_w_0_s1_writedata),     //                                                           .writedata
		.data_tx_to_w_0_s1_chipselect                                     (mm_interconnect_0_data_tx_to_w_0_s1_chipselect),    //                                                           .chipselect
		.fsm_info_s1_address                                              (mm_interconnect_0_fsm_info_s1_address),             //                                                fsm_info_s1.address
		.fsm_info_s1_readdata                                             (mm_interconnect_0_fsm_info_s1_readdata),            //                                                           .readdata
		.fsm_info_0_s1_address                                            (mm_interconnect_0_fsm_info_0_s1_address),           //                                              fsm_info_0_s1.address
		.fsm_info_0_s1_readdata                                           (mm_interconnect_0_fsm_info_0_s1_readdata),          //                                                           .readdata
		.led_fpga_s1_address                                              (mm_interconnect_0_led_fpga_s1_address),             //                                                led_fpga_s1.address
		.led_fpga_s1_write                                                (mm_interconnect_0_led_fpga_s1_write),               //                                                           .write
		.led_fpga_s1_readdata                                             (mm_interconnect_0_led_fpga_s1_readdata),            //                                                           .readdata
		.led_fpga_s1_writedata                                            (mm_interconnect_0_led_fpga_s1_writedata),           //                                                           .writedata
		.led_fpga_s1_chipselect                                           (mm_interconnect_0_led_fpga_s1_chipselect),          //                                                           .chipselect
		.link_disable_s1_address                                          (mm_interconnect_0_link_disable_s1_address),         //                                            link_disable_s1.address
		.link_disable_s1_write                                            (mm_interconnect_0_link_disable_s1_write),           //                                                           .write
		.link_disable_s1_readdata                                         (mm_interconnect_0_link_disable_s1_readdata),        //                                                           .readdata
		.link_disable_s1_writedata                                        (mm_interconnect_0_link_disable_s1_writedata),       //                                                           .writedata
		.link_disable_s1_chipselect                                       (mm_interconnect_0_link_disable_s1_chipselect),      //                                                           .chipselect
		.link_disable_0_s1_address                                        (mm_interconnect_0_link_disable_0_s1_address),       //                                          link_disable_0_s1.address
		.link_disable_0_s1_write                                          (mm_interconnect_0_link_disable_0_s1_write),         //                                                           .write
		.link_disable_0_s1_readdata                                       (mm_interconnect_0_link_disable_0_s1_readdata),      //                                                           .readdata
		.link_disable_0_s1_writedata                                      (mm_interconnect_0_link_disable_0_s1_writedata),     //                                                           .writedata
		.link_disable_0_s1_chipselect                                     (mm_interconnect_0_link_disable_0_s1_chipselect),    //                                                           .chipselect
		.link_start_s1_address                                            (mm_interconnect_0_link_start_s1_address),           //                                              link_start_s1.address
		.link_start_s1_write                                              (mm_interconnect_0_link_start_s1_write),             //                                                           .write
		.link_start_s1_readdata                                           (mm_interconnect_0_link_start_s1_readdata),          //                                                           .readdata
		.link_start_s1_writedata                                          (mm_interconnect_0_link_start_s1_writedata),         //                                                           .writedata
		.link_start_s1_chipselect                                         (mm_interconnect_0_link_start_s1_chipselect),        //                                                           .chipselect
		.link_start_0_s1_address                                          (mm_interconnect_0_link_start_0_s1_address),         //                                            link_start_0_s1.address
		.link_start_0_s1_write                                            (mm_interconnect_0_link_start_0_s1_write),           //                                                           .write
		.link_start_0_s1_readdata                                         (mm_interconnect_0_link_start_0_s1_readdata),        //                                                           .readdata
		.link_start_0_s1_writedata                                        (mm_interconnect_0_link_start_0_s1_writedata),       //                                                           .writedata
		.link_start_0_s1_chipselect                                       (mm_interconnect_0_link_start_0_s1_chipselect),      //                                                           .chipselect
		.MONITOR_A_s1_address                                             (mm_interconnect_0_monitor_a_s1_address),            //                                               MONITOR_A_s1.address
		.MONITOR_A_s1_readdata                                            (mm_interconnect_0_monitor_a_s1_readdata),           //                                                           .readdata
		.MONITOR_B_s1_address                                             (mm_interconnect_0_monitor_b_s1_address),            //                                               MONITOR_B_s1.address
		.MONITOR_B_s1_readdata                                            (mm_interconnect_0_monitor_b_s1_readdata),           //                                                           .readdata
		.send_fct_now_s1_address                                          (mm_interconnect_0_send_fct_now_s1_address),         //                                            send_fct_now_s1.address
		.send_fct_now_s1_write                                            (mm_interconnect_0_send_fct_now_s1_write),           //                                                           .write
		.send_fct_now_s1_readdata                                         (mm_interconnect_0_send_fct_now_s1_readdata),        //                                                           .readdata
		.send_fct_now_s1_writedata                                        (mm_interconnect_0_send_fct_now_s1_writedata),       //                                                           .writedata
		.send_fct_now_s1_chipselect                                       (mm_interconnect_0_send_fct_now_s1_chipselect),      //                                                           .chipselect
		.send_fct_now_0_s1_address                                        (mm_interconnect_0_send_fct_now_0_s1_address),       //                                          send_fct_now_0_s1.address
		.send_fct_now_0_s1_write                                          (mm_interconnect_0_send_fct_now_0_s1_write),         //                                                           .write
		.send_fct_now_0_s1_readdata                                       (mm_interconnect_0_send_fct_now_0_s1_readdata),      //                                                           .readdata
		.send_fct_now_0_s1_writedata                                      (mm_interconnect_0_send_fct_now_0_s1_writedata),     //                                                           .writedata
		.send_fct_now_0_s1_chipselect                                     (mm_interconnect_0_send_fct_now_0_s1_chipselect),    //                                                           .chipselect
		.timec_en_to_tx_s1_address                                        (mm_interconnect_0_timec_en_to_tx_s1_address),       //                                          timec_en_to_tx_s1.address
		.timec_en_to_tx_s1_write                                          (mm_interconnect_0_timec_en_to_tx_s1_write),         //                                                           .write
		.timec_en_to_tx_s1_readdata                                       (mm_interconnect_0_timec_en_to_tx_s1_readdata),      //                                                           .readdata
		.timec_en_to_tx_s1_writedata                                      (mm_interconnect_0_timec_en_to_tx_s1_writedata),     //                                                           .writedata
		.timec_en_to_tx_s1_chipselect                                     (mm_interconnect_0_timec_en_to_tx_s1_chipselect),    //                                                           .chipselect
		.timec_en_to_tx_0_s1_address                                      (mm_interconnect_0_timec_en_to_tx_0_s1_address),     //                                        timec_en_to_tx_0_s1.address
		.timec_en_to_tx_0_s1_write                                        (mm_interconnect_0_timec_en_to_tx_0_s1_write),       //                                                           .write
		.timec_en_to_tx_0_s1_readdata                                     (mm_interconnect_0_timec_en_to_tx_0_s1_readdata),    //                                                           .readdata
		.timec_en_to_tx_0_s1_writedata                                    (mm_interconnect_0_timec_en_to_tx_0_s1_writedata),   //                                                           .writedata
		.timec_en_to_tx_0_s1_chipselect                                   (mm_interconnect_0_timec_en_to_tx_0_s1_chipselect),  //                                                           .chipselect
		.timec_rx_r_s1_address                                            (mm_interconnect_0_timec_rx_r_s1_address),           //                                              timec_rx_r_s1.address
		.timec_rx_r_s1_readdata                                           (mm_interconnect_0_timec_rx_r_s1_readdata),          //                                                           .readdata
		.timec_rx_r_0_s1_address                                          (mm_interconnect_0_timec_rx_r_0_s1_address),         //                                            timec_rx_r_0_s1.address
		.timec_rx_r_0_s1_readdata                                         (mm_interconnect_0_timec_rx_r_0_s1_readdata),        //                                                           .readdata
		.timec_rx_ready_s1_address                                        (mm_interconnect_0_timec_rx_ready_s1_address),       //                                          timec_rx_ready_s1.address
		.timec_rx_ready_s1_readdata                                       (mm_interconnect_0_timec_rx_ready_s1_readdata),      //                                                           .readdata
		.timec_rx_ready_0_s1_address                                      (mm_interconnect_0_timec_rx_ready_0_s1_address),     //                                        timec_rx_ready_0_s1.address
		.timec_rx_ready_0_s1_readdata                                     (mm_interconnect_0_timec_rx_ready_0_s1_readdata),    //                                                           .readdata
		.timec_tx_ready_s1_address                                        (mm_interconnect_0_timec_tx_ready_s1_address),       //                                          timec_tx_ready_s1.address
		.timec_tx_ready_s1_readdata                                       (mm_interconnect_0_timec_tx_ready_s1_readdata),      //                                                           .readdata
		.timec_tx_ready_0_s1_address                                      (mm_interconnect_0_timec_tx_ready_0_s1_address),     //                                        timec_tx_ready_0_s1.address
		.timec_tx_ready_0_s1_readdata                                     (mm_interconnect_0_timec_tx_ready_0_s1_readdata),    //                                                           .readdata
		.timec_tx_to_w_s1_address                                         (mm_interconnect_0_timec_tx_to_w_s1_address),        //                                           timec_tx_to_w_s1.address
		.timec_tx_to_w_s1_write                                           (mm_interconnect_0_timec_tx_to_w_s1_write),          //                                                           .write
		.timec_tx_to_w_s1_readdata                                        (mm_interconnect_0_timec_tx_to_w_s1_readdata),       //                                                           .readdata
		.timec_tx_to_w_s1_writedata                                       (mm_interconnect_0_timec_tx_to_w_s1_writedata),      //                                                           .writedata
		.timec_tx_to_w_s1_chipselect                                      (mm_interconnect_0_timec_tx_to_w_s1_chipselect),     //                                                           .chipselect
		.timec_tx_to_w_0_s1_address                                       (mm_interconnect_0_timec_tx_to_w_0_s1_address),      //                                         timec_tx_to_w_0_s1.address
		.timec_tx_to_w_0_s1_write                                         (mm_interconnect_0_timec_tx_to_w_0_s1_write),        //                                                           .write
		.timec_tx_to_w_0_s1_readdata                                      (mm_interconnect_0_timec_tx_to_w_0_s1_readdata),     //                                                           .readdata
		.timec_tx_to_w_0_s1_writedata                                     (mm_interconnect_0_timec_tx_to_w_0_s1_writedata),    //                                                           .writedata
		.timec_tx_to_w_0_s1_chipselect                                    (mm_interconnect_0_timec_tx_to_w_0_s1_chipselect)    //                                                           .chipselect
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~hps_0_h2f_reset_reset),             // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
